User|Original_User/Web|Compound|Negative|Neutral|Positive|Tweet
GoldenbergLaw|twinsational|-0.0258|0.136|0.734|0.13|RT @twinsational: A #Trump Fan Just Pulled A Gun On A Black Voter At #Florida Polling Station - https://t.co/fstiatqr1o
GoldenbergLaw|occupydemocrats|-0.0258|0.136|0.734|0.13|RT @twinsational: A #Trump Fan Just Pulled A Gun On A Black Voter At #Florida Polling Station - https://t.co/fstiatqr1o
MachPierogi|syoka68|-0.2462|0.099|0.901|0.0|RT @syoka68: Not hard to believe they are rigging exit polls! Turn off the tv GO VOTE TRUMP! https://t.co/HLNXmSp0IQ
MachPierogi|twitter|-0.2462|0.099|0.901|0.0|RT @syoka68: Not hard to believe they are rigging exit polls! Turn off the tv GO VOTE TRUMP! https://t.co/HLNXmSp0IQ
GodlessNZ|itsugamom|0.6093|0.0|0.819|0.181|RT @itsugamom: #StayInLine ....So proud of Trumpsters! Just take a fold out chair! When you vote Trump we will #DrainTheSwamp! 
iAmsterdamNews|christianitytoday|0.2023|0.0|0.878|0.122|Top 10 Stats Explaining the Evangelical Vote for Trump or Clinton https://t.co/iRbj1bZRjw #Amsterdam #News
NJbyMarriage|NivenJ1|-0.9001|0.5|0.5|0.0|RT @NivenJ1: Trump: I hate illegal immigrants.Melania: 'I hate cyber bullies'*look at each other longingly*
jamesfoxx19|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
Artco77|guitarboyjohnny|0.0|0.0|1.0|0.0|RT @guitarboyjohnny: Trump leads Clinton 32 to 25 votes in New Hampshire. EVERYONE TO CANADA!!!
Morwennnnna|TheLadBible|0.3612|0.0|0.848|0.152|RT @TheLadBible: Stevie Wonder says Trump being President is like him driving a car. https://t.co/cpaF7yRJdz https://t.co/WcW5NvNcWv
Morwennnnna|theladbible|0.3612|0.0|0.848|0.152|RT @TheLadBible: Stevie Wonder says Trump being President is like him driving a car. https://t.co/cpaF7yRJdz https://t.co/WcW5NvNcWv
mythicalbellamy|BlakeBeMine|-0.6486|0.389|0.474|0.137|RT @BlakeBeMine: Accuse me of supporting Trump and I'll block your ass so fast
bitterflie|pattonoswalt|0.0|0.0|1.0|0.0|RT @pattonoswalt: OMG Donald Trump just texted this to me. Does he already know I voted for Clinton? https://t.co/7COBWg7imR
bitterflie|twitter|0.0|0.0|1.0|0.0|RT @pattonoswalt: OMG Donald Trump just texted this to me. Does he already know I voted for Clinton? https://t.co/7COBWg7imR
WhittyWhit86|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
WhittyWhit86|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
EchoesOfKyraaa|Big_Shug99|0.8316|0.0|0.729|0.271|RT @Big_Shug99: So is there an application for head cotton picker if Trump wins. I think I have great management skills to get cotton picke
philboldt|NoahCRothman|-0.1531|0.157|0.714|0.129|@NoahCRothman @BanditGolf @NewsPolitics Maybe if Trump would of insulted a few more people. That could of help right?
MGlick78|BillGalston|0.5859|0.0|0.847|0.153|"RT @BillGalston: Early exit polls show Trump and Clinton are neck-and-neck among whites with a college degree. If Dems win this group, hist"
sirdrano|livelrod|0.0|0.0|1.0|0.0|RT @livelrod: Voted! #TRUMP https://t.co/09MmBBVWYg
sirdrano|twitter|0.0|0.0|1.0|0.0|RT @livelrod: Voted! #TRUMP https://t.co/09MmBBVWYg
tamaraleighllc|trfgrp|0.0|0.0|1.0|0.0|"RT @trfgrp: Our projection: Trump 306 Clinton 223 w/CO, VA &amp; WI possibly breaking Trump as ""hidden voter"" #trumptiderolls https://t.co/u34D"
tamaraleighllc|t|0.0|0.0|1.0|0.0|"RT @trfgrp: Our projection: Trump 306 Clinton 223 w/CO, VA &amp; WI possibly breaking Trump as ""hidden voter"" #trumptiderolls https://t.co/u34D"
Larkell_|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
fredbauerblog|nationalreview|0.0|0.0|1.0|0.0|"Before the deluge of results, I'll reiterate this: Our republic will survive whatever the result. https://t.co/TUW7beveWb"
election_votes|C_Smatana|0.0|0.0|1.0|0.0|RT @C_Smatana: Who are you voting for Trump or Clinton?!? #ElectionDay #USElection2016 #ElectionNight #HillaryClintonForPresident #DonaldTr
mottstreet6|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
thatdaba|TheLastRefuge2|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
thatdaba|twitter|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
clodma0202|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
stratocat1012|Bikers4Trump|-0.6486|0.227|0.773|0.0|RT @Bikers4Trump: We need Trump &amp; #ImVotingBecause @HillaryClinton is a criminal &amp; must be stopped this Election Eve#RETWEET &amp; Visit https
nutifafa_max|Ryan23675317|0.4767|0.098|0.675|0.227|RT @Ryan23675317: Just in case trump wins I'm latin btw I'll miss yall
rhinoceroseosei|Bill_Nye_Tho|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
rhinoceroseosei|twitter|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
johnboor|BillMoyers|0.0|0.0|1.0|0.0|Trumps Three Biggest Enablers - https://t.co/HnJY9Rgfnp https://t.co/QywMDcYgks
boredhoney|SteadyTheo|0.4939|0.0|0.868|0.132|"RT @SteadyTheo: Drink water, don't vote for Donald Trump, express empathy, enjoy art,  don't compare yourself to other people, do not read"
FranP20|nytpolitics|-0.7783|0.302|0.698|0.0|@nytpolitics ppl say that Trump plans a class action lawsuit against anyone who did not vote for him. He's just a Sore Loser.
TheoJans1|MMFlint|0.05|0.105|0.782|0.113|Hear hear @MMFlint Do vote dear Americans. But not for #Trump Thanks on behalf of the people of the Netherlands.
Deibliane1|mitchellvii|0.0|0.0|1.0|0.0|@mitchellvii this County is heavy for Trump
mkearley2008|WardahHashmi|0.0|0.0|1.0|0.0|@WardahHashmi Look who's she's running against. I don't think Trump could find Pakistan on a map.
sherrymisner|dawg_lb|0.0|0.0|1.0|0.0|"RT @dawg_lb: Hillary R Clinton,YOU SHOULD NEVER BE ABLE TO LOOK AT YOURSELF IN THE MIRROR!!!!!!!VOTE AS FAST AS YOU CAN!!!!!!!!!!TRUM"
torres_dalkin|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
torres_dalkin|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
Pell48|RosieBud521|0.3296|0.214|0.614|0.172|RT @RosieBud521: No @MegynKelly tonight!  I can't stand her hatred and bias against Trump! @SeanHannity https://t.co/4QJC1ll74U
Pell48|twitter|0.3296|0.214|0.614|0.172|RT @RosieBud521: No @MegynKelly tonight!  I can't stand her hatred and bias against Trump! @SeanHannity https://t.co/4QJC1ll74U
truenorth_eh|tamaraleighllc|0.4019|0.0|0.828|0.172|RT @tamaraleighllc: Yes I did  VOTED #Trump  #ElectionDay #WI #Wisconsin #MAGA #NeverHillary @AmericaFirst #DrainTheSwamp #WomenForT
mr_burton23|RawStory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
mr_burton23|rawstory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
louulevv1|evrydayfeminism|0.5994|0.0|0.671|0.329|Dear White America: You Are All Responsible for Trump https://t.co/39y18LV26z via @evrydayfeminism
louulevv1|everydayfeminism|0.5994|0.0|0.671|0.329|Dear White America: You Are All Responsible for Trump https://t.co/39y18LV26z via @evrydayfeminism
nicholas51|newsmax|0.0|0.0|1.0|0.0|"RT @newsmax: With 1% of the vote in for Kentucky, Trump is holding a steady lead over Hillary Clinton. #ElectionNight #myvote2016 https://t"
nicholas51||0.0|0.0|1.0|0.0|"RT @newsmax: With 1% of the vote in for Kentucky, Trump is holding a steady lead over Hillary Clinton. #ElectionNight #myvote2016 https://t"
cmrose999|VoteStand|0.0|0.0|1.0|0.0|"RT @VoteStand: Tucson, AZ: ""Tucson poll workers telling a Hispanic woman (my wife) that she would be deported if she voted for Trump."""
myecoll|NaYaKnoMi|-0.1779|0.086|0.914|0.0|"RT @NaYaKnoMi: i can't believe people are actually voting for trump. seriously, it is happening... they're voting for a clinically certifie"
tlynn561|kayleighmcenany|0.0|0.0|1.0|0.0|RT @kayleighmcenany: Evening voters could determine this election - you still have time to go vote Trump!!!  #ElectionNight
WilliamSDraper|JRehling|0.4939|0.08|0.725|0.196|RT @JRehling: When is Obama supposed to take everyone's guns and impose Islamic law? The people supporting Trump now promised us that 4 and
feltonewt|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
lilaustin110|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
blurrygambino|twitter|0.128|0.169|0.635|0.196|When you realize that we're screwed if trump or Hillary wins the election https://t.co/5ULRBFJVIR
courtalexandra_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
punksandwitch|bernorjill|0.707|0.124|0.473|0.402|"RT @bernorjill: Dear Clinton Supporter, I Don't Care If You're Afraid Of A Trump Win https://t.co/GVmxpbqkEF"
punksandwitch|progressivearmy|0.707|0.124|0.473|0.402|"RT @bernorjill: Dear Clinton Supporter, I Don't Care If You're Afraid Of A Trump Win https://t.co/GVmxpbqkEF"
Activeviii|FrankLuntz|-0.1027|0.055|0.945|0.0|RT @FrankLuntz: The turnout in Democratic Philadelphia is so high that it's hard to see Trump overcoming it in the rest of the state.  #Ele
welzZalia|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
CiroacardenasA|nytimes|0.1098|0.177|0.633|0.19|"RT @nytimes: ""If we don't win, this will be the single greatest waste of time, energy and money in my life,"" Donald Trump said https://t.co"
CiroacardenasA|t|0.1098|0.177|0.633|0.19|"RT @nytimes: ""If we don't win, this will be the single greatest waste of time, energy and money in my life,"" Donald Trump said https://t.co"
steve2blue4u|JaredWyand|0.8481|0.0|0.495|0.505|@JaredWyand not a New England or Brady fan but glad 2 c them support Trump
BBCARKING|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
ColdestCorazon|MostDopeSince94|0.0772|0.0|0.915|0.085|RT @MostDopeSince94: i don't understand how you can be a minority n still want to vote for trump...
sargentolipton|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
hlewissss|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
chelseajae1103|jcrum417|0.2023|0.0|0.921|0.079|@jcrum417 @AffinityxD @DrJillStein the elite are the people in power. Both government and market. And Hilary and trump are playing both side
NoelleTMD|trump_woman|0.4199|0.0|0.787|0.213|RT @trump_woman: 10-Foot-Tall TRUMP! Letters Greet Los Angeles Highway 101 Freeway Commuters https://t.co/0OZz0U1vpb via @trump_woman #Ca
NoelleTMD|losangeles|0.4199|0.0|0.787|0.213|RT @trump_woman: 10-Foot-Tall TRUMP! Letters Greet Los Angeles Highway 101 Freeway Commuters https://t.co/0OZz0U1vpb via @trump_woman #Ca
lonireeder|ClaireB20164206|0.0|0.0|1.0|0.0|@ClaireB20164206 Trump voters believe they'll all get a new doublewide &amp; a case of beer if they vote 4 him! (remodeled outhouses too!) 
AveEuropa|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
AveEuropa|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
JehseaLynn|JuddLegum|-0.1027|0.128|0.765|0.107|RT @JuddLegum: Trump black outreach strategy:1. Your lives are miserable2. You have nothing to lose3. Beyonc sucks
skorpyos|TeaPartyCat|-0.547|0.22|0.714|0.066|"RT @TeaPartyCat: It's not fair to call all Trump's supporters racist and sexist. Some are racist, some are sexist, but not all of them are"
dr3am_ch4sing|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
dr3am_ch4sing|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Zackdjohnson1|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
Zackdjohnson1|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
tashaaamay|LouisePentland|0.4926|0.0|0.856|0.144|"RT @LouisePentland: Going to bed. When I wake up, Trump better not be the President or I'm going back to sleep!"
FosterNeegreen|pchowder|-0.7506|0.262|0.738|0.0|RT @pchowder: understand why #Trump is pissed off at #GOP-drove past NHGOP headquarters a dozen people holding #KellyAyotte signs- no one e
StarmanRock|LouDobbs|0.6249|0.0|0.683|0.317|@LouDobbs @kimguilfoyle @EdRollins @mgoodwin_nypost @tony4ny @lh_carter will do. We want watch Trump win
mental_nigella_|discokidnap|0.0|0.0|1.0|0.0|RT @discokidnap: Bet Sunderland votes for Trump.
riddlepots|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
riddlepots|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
nordicscripts|hrtablaze|0.5399|0.0|0.868|0.132|RT @hrtablaze: CNN reporting that there is record breaking turnout! That is good news for the Trump Train ! First Exit Poll comes out short
TherealMelHall|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
prairiepoultry|CBSEveningNews|0.6705|0.0|0.766|0.234|"@CBSEveningNews  Nice job of portraying only Trump as the ""deplorable"" candidate in your special. Clinton deserves some of that ""limelight """
DrThomasPaul|DrThomasPaul|-0.1531|0.164|0.701|0.136|"RT @DrThomasPaul: .@HillarysAmerica is one of division, crime, #pharma &amp; riots.It's good for corrupt #BigBusiness.#gmo #Hillary #Trumphttp"
JohnRCurtis|LordAshcroft|0.0|0.0|1.0|0.0|RT @LordAshcroft: Early US exit polls. Georgia Trump +3. Virginia Clinton+8. N. Carolina Clinton+2. Ohio Tie. Florida Clinton +2. New Hamps
Friday_Everyday|CryingJordan|0.0|0.0|1.0|0.0|RT @CryingJordan: A Donald Trump cake being wheeled into Trump Tower #ElectionDay https://t.co/9kVYIKgZ5d
Friday_Everyday|twitter|0.0|0.0|1.0|0.0|RT @CryingJordan: A Donald Trump cake being wheeled into Trump Tower #ElectionDay https://t.co/9kVYIKgZ5d
enfingercolton2|mitchellvii|0.4404|0.0|0.805|0.195|"RT @mitchellvii: Trump leads IND 72-25.  Good Lord people, something is happening here."
BeatsBy777|UglyGod|-0.5106|0.121|0.879|0.0|RT @UglyGod: It means yall shoulda fuckin listened &amp; kept Bernie Sanders as an option cause now we all look dumb af choosing between Hillar
lwtsheeran|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
McMystie|twitter|0.0|0.0|1.0|0.0|#FoxNews2016 #Election2016 #MAGA Our 6 year old voted Trump! https://t.co/Y1TOR9Cr3v
LVJudy89128|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Maddman1212|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
Maddman1212|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
jbisrael|igorbobic|-0.4588|0.167|0.833|0.0|"RT @igorbobic: NV judge calls Trump campaign request to preserve poll data in Clark County offensive"""
Sublyminal12|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
celiaj02|GartrellLinda|0.2714|0.0|0.905|0.095|RT @GartrellLinda: Important! RTGET OUT THERE &amp; VOTE TRUMPSTERSVERY TIGHT in Florida panhandle. Call everyone you know to get those Trump
rapidcraft|realDonaldTrump|-0.4215|0.219|0.781|0.0|"Report: Voter Intimidation in Philly, @realDonaldTrump Observers Kicked Out https://t.co/jqoZLU0INP @Phillydotcom"
rapidcraft|infowars|-0.4215|0.219|0.781|0.0|"Report: Voter Intimidation in Philly, @realDonaldTrump Observers Kicked Out https://t.co/jqoZLU0INP @Phillydotcom"
sheacollagen|uniqueprophet|0.0258|0.153|0.691|0.157|"RT @uniqueprophet: OOPS @realDonaldTrump, @trump TRUMP SUPPORTERS, WE HAVE ENDURED TOO MUCH STRESS, EMOTION,EFFORT,DON'T LET LEFT SCUM STEA"
APOYODECHILE|mitchellvii|0.2177|0.137|0.684|0.179|RT @mitchellvii: So was Trump winning CO and conveniently every voting machine in the state broke?
cowboycoffee|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
cowboycoffee|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
ruthe_susan|Wil_Johnson1|0.0|0.0|1.0|0.0|"RT @Wil_Johnson1: In Kentucky and Indiana with just a little over 3% reporting, Trump is getting 2-1 votes over Hillary https://t.co/4wCD0Q"
ruthe_susan|t|0.0|0.0|1.0|0.0|"RT @Wil_Johnson1: In Kentucky and Indiana with just a little over 3% reporting, Trump is getting 2-1 votes over Hillary https://t.co/4wCD0Q"
cnsltngmexican|Bill_Nye_Tho|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
cnsltngmexican|twitter|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
BurrRobson|Trump_Videos|-0.5423|0.22|0.78|0.0|@Trump_Videos No loss in my opinion. She should have been born in the USSR and headed the KGB.
OneLoveManUtd|Deadspin|0.0|0.0|1.0|0.0|RT @Deadspin: The Trump campaign wants to make names of Nevada poll workers public. Judge's response: https://t.co/tes99IMbbH
OneLoveManUtd|twitter|0.0|0.0|1.0|0.0|RT @Deadspin: The Trump campaign wants to make names of Nevada poll workers public. Judge's response: https://t.co/tes99IMbbH
atf13atf|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Cheddabob101|RubenAbeyta|-0.8625|0.591|0.303|0.106|"@RubenAbeyta no you offended me Fuck you, you racist trump supporter"
TwinParasite|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
TwinParasite|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
bIanceclare|pearlwillam|0.4404|0.0|0.847|0.153|RT @pearlwillam: @CeeJayCraig i would've aborted them if i knew they were gonna grow up to be trump supporters
billybudd16|renata_piranha|-0.7339|0.27|0.73|0.0|RT @renata_piranha: @jornalnacional @realDonaldTrump  BREAKING:MachineRefuses toAllow VoteFor Trump in Pennsylvania!!RT the hell out of it
Lydon93|BtheHill|0.4588|0.115|0.673|0.212|"RT @BtheHill: I hope if Trump wins his first words of his inaugural speech are going to be ""You're Fired"" with a finger pointed directly at"
keluttcu|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
dougsmith1946|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
JoCastiglione|Trumpocrats|0.0|0.0|1.0|0.0|RT @Trumpocrats: Reuters showing a surge #ElectionDay #ElectionNight #DrainTheSwamp #MAGA3X #LANDSLIDE #PodestaEmails #Trump https://t.co/A
JoCastiglione|amandeep|0.0|0.0|1.0|0.0|RT @Trumpocrats: Reuters showing a surge #ElectionDay #ElectionNight #DrainTheSwamp #MAGA3X #LANDSLIDE #PodestaEmails #Trump https://t.co/A
katherinems00|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
katherinems00|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
natalieeeemary|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
bmcpa85|GovMikeHuckabee|-0.0516|0.059|0.941|0.0|"RT @GovMikeHuckabee: I personally know both candidates;Have for years; Not hard choice. Neither are perfect-nor am I, but voted Trump w/o h"
KennethClayden|LukeIsNotSexy|0.25|0.0|0.92|0.08|"@LukeIsNotSexy Not the time for jokes, Luke, we could be looking at a Trump presidency if a few people (I don't know the actual figure) did"
TonyTalbo|oreillyfactor|0.0|0.0|1.0|0.0|Rigging #176 Broward #RiggedSystem #TRUMP #TrumpPence16 #draintheswamp #MAGA #TrumpTrain @oreillyfactor https://t.co/e4nsdBlWMq
TonyTalbo|twitter|0.0|0.0|1.0|0.0|Rigging #176 Broward #RiggedSystem #TRUMP #TrumpPence16 #draintheswamp #MAGA #TrumpTrain @oreillyfactor https://t.co/e4nsdBlWMq
AnonBruja|nealrogers|-0.4981|0.123|0.877|0.0|RT @nealrogers: Trump says Tom Brady told him hed voted for him. Brady says he hasnt voted yet; wife Gisele Bundchen answers NO! https:
MonaBuckmiller|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
MonaBuckmiller|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
Teressastone4|joelpollak|0.4019|0.0|0.838|0.162|RT @joelpollak: Trump Fans Sing Star-Spangled Banner in Front of Victory Party https://t.co/wVlNFT9hzp via @BreitbartNews
Teressastone4|breitbart|0.4019|0.0|0.838|0.162|RT @joelpollak: Trump Fans Sing Star-Spangled Banner in Front of Victory Party https://t.co/wVlNFT9hzp via @BreitbartNews
dangstephen2sa1|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
dangstephen2sa1|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
Tutoanana|SteveRattner|-0.0258|0.152|0.702|0.146|RT @SteveRattner: Exit polls: border wall54% oppose 40% supportLooks like a losing issue for Trump#Election2016
F_kFlyImFashion|Iemonade|0.3939|0.0|0.84|0.16|"RT @Iemonade: trump voters in the hive ?? come up to the mic, please. https://t.co/AuT29iQLe2"
F_kFlyImFashion|twitter|0.3939|0.0|0.84|0.16|"RT @Iemonade: trump voters in the hive ?? come up to the mic, please. https://t.co/AuT29iQLe2"
tabykinz|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
MarioHazelwood|ZachAJacobson|0.8625|0.0|0.676|0.324|"RT @ZachAJacobson: Yes, I voted Hillary. You voted Trump? Nice. Won't change how I, or anybody else should view you. Great thing about Amer"
OneTrump4All|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
OneTrump4All|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
LESTERHICKEYS|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
LESTERHICKEYS|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
kLodeserto|mitchellvii|0.2177|0.137|0.684|0.179|RT @mitchellvii: So was Trump winning CO and conveniently every voting machine in the state broke?
naezzy_|heartless_haze|-0.1027|0.195|0.632|0.172|RT @heartless_haze: Whoever voted for Trump is honestly as stupid as he is
UnitedBrews|EireKav|0.0|0.0|1.0|0.0|RT @EireKav: Kentucky get out and VOTE Trump. This might be BS to make you believe its in the bag. It is NOT until everyone who can votes f
SergiosWisdom|AmericasVoice|-0.2023|0.094|0.848|0.058|RT @AmericasVoice: BREAKING: National exit poll number for Latino Voters from @LatinoDecisions: Clinton 79 - Trump 18. New low for GOP. Sam
Jakelopz17|CBSNews|0.0|0.0|1.0|0.0|"RT @CBSNews: If Donald Trump were elected, this is how he would impact your taxes. https://t.co/T49gkrVAlv"
Jakelopz17|twitter|0.0|0.0|1.0|0.0|"RT @CBSNews: If Donald Trump were elected, this is how he would impact your taxes. https://t.co/T49gkrVAlv"
1blessedbee|healthandcents|-0.41|0.215|0.671|0.113|"RT @healthandcents: @payao1a1 ABSOLUTE TRUTH. If #Trump does not win this, we will never have free election again. #Globalists will control"
AshtonLigan|KayleePages|0.5499|0.0|0.785|0.215|"@KayleePages but many wish trump can just be shot already, it was already attempted"
RHYDOE|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
RHYDOE|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Cricaholics|itvnews|0.0|0.0|1.0|0.0|RT @itvnews: US Election: Stark difference between how men and women are expected to vote #Election2016 #ElectionNight https://t.co/BfQPcj2
Cricaholics|t|0.0|0.0|1.0|0.0|RT @itvnews: US Election: Stark difference between how men and women are expected to vote #Election2016 #ElectionNight https://t.co/BfQPcj2
EmilVelour|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
mwarhurst|DenisMacShane|-0.2263|0.153|0.766|0.08|RT @DenisMacShane: Quelle surprise. Unlike the Leave Lies in Brexit unchallenged by BBC and transmitted by most press Trump has not been gi
LiberalRevival|businessinsider|0.0|0.0|1.0|0.0|RT @businessinsider: Donald Trumps outlandish persona might be due to his decades-long relationship with @WWE #ElectionNight https://t.c
LiberalRevival||0.0|0.0|1.0|0.0|RT @businessinsider: Donald Trumps outlandish persona might be due to his decades-long relationship with @WWE #ElectionNight https://t.c
elitetech333|LarrySchweikart|0.0|0.0|1.0|0.0|"@LarrySchweikart my 5 CO-workers and their spouses, ALL TRUMP!!!"
angela_rose06|JYSexton|-0.5975|0.175|0.825|0.0|"RT @JYSexton: Donald Trump and the forces of bigotry are counting on you not caring, on you not exercising your rights, on you not trusting"
Liana_Guerra|MarcACaputo|-0.1531|0.138|0.748|0.114|RT @MarcACaputo: Good news for Clinton and ergo bad news for Trump in FL's most Democratic performing major urban county https://t.co/L3qZv
Liana_Guerra|t|-0.1531|0.138|0.748|0.114|RT @MarcACaputo: Good news for Clinton and ergo bad news for Trump in FL's most Democratic performing major urban county https://t.co/L3qZv
maweypooh1|JaredWyand|-0.5574|0.167|0.833|0.0|RT @JaredWyand: She's caught paying people to riot at Trump ralliesHer whole inner circle does Satanic #SpiritCookingAnd last night...
Anaruiz415|litzymarie_|0.8225|0.0|0.648|0.352|"RT @litzymarie_: if trump wins today, im taking myself to mexico even tho i got papers lmao"
Kencarterpounds|HillaryClinton|0.296|0.223|0.446|0.33|"@HillaryClinton You have won, Trump is a mess"
itunes65|mitchellvii|0.5267|0.0|0.673|0.327|RT @mitchellvii: I see Trump winning MI and CO.
BusinessNews40|businessinsider|0.4588|0.117|0.612|0.27|"Donald Trump's website was saying some odd things, thanks to a security hole https://t.co/2IeBqY1DyX #Business https://t.co/Fag5u71SCg"
swaggiemario|yuppjulian|0.4648|0.0|0.822|0.178|RT @yuppjulian: BEFORE TRUMP BECOMES PRESIDENT MAKE SURE YOU WATCH MY NEW VIDEO https://t.co/Bdtz0KP3Hl #goonsnewvideo
swaggiemario|youtube|0.4648|0.0|0.822|0.178|RT @yuppjulian: BEFORE TRUMP BECOMES PRESIDENT MAKE SURE YOU WATCH MY NEW VIDEO https://t.co/Bdtz0KP3Hl #goonsnewvideo
kianajones200|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
kianajones200|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
dcas1978|AmericasVoice|-0.2023|0.094|0.848|0.058|RT @AmericasVoice: BREAKING: National exit poll number for Latino Voters from @LatinoDecisions: Clinton 79 - Trump 18. New low for GOP. Sam
lblink949|lisserlou47|0.5719|0.0|0.856|0.144|"RT @lisserlou47: @DonaldJTrumpJr when I voted TRUMP I did not vote for dem or rep, I voted for a MAN that loves America and has given and s"
JimmyJames38|nbc4i|0.0|0.0|1.0|0.0|RT @nbc4i: 102-year-old woman casts her vote for Donald Trump. https://t.co/rhJNJSy0rf https://t.co/jmz9hMN9YY
JimmyJames38|nbc4i|0.0|0.0|1.0|0.0|RT @nbc4i: 102-year-old woman casts her vote for Donald Trump. https://t.co/rhJNJSy0rf https://t.co/jmz9hMN9YY
gdg2024|mitchellvii|0.4404|0.0|0.838|0.162|"RT @mitchellvii: If Trump ends up dramatically outperfroming his RCP averages in early states, good sign."
mmcandy64|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
KashItIs|twitter|0.128|0.0|0.88|0.12|"It's on your snap, everyone knows you voted Trump you supremacist https://t.co/t10fzyv1kb"
Mikehall73|RealJamesWoods|0.5411|0.0|0.696|0.304|@RealJamesWoods In honor of you Mr Woods.  Trump! https://t.co/OKMTgDd8dE
Mikehall73|twitter|0.5411|0.0|0.696|0.304|@RealJamesWoods In honor of you Mr Woods.  Trump! https://t.co/OKMTgDd8dE
NRodibaugh|mmfafa|0.5267|0.103|0.647|0.25|"RT @mmfafa: Fox News just played the ""Blame Russia"" Card...Trump MUST be winning. @mitchellvii @Cernovich @AwesomeIva @StefanMolyneux @Pris"
trapgod_Ben|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
trapgod_Ben|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
boogeyone|Scout_Finch|0.0258|0.156|0.684|0.16|RT @Scout_Finch: I will remember you. Will you remember me? In memoriam ... the best of the worst Trump pundits https://t.co/J04tJ28yfG
boogeyone|twitter|0.0258|0.156|0.684|0.16|RT @Scout_Finch: I will remember you. Will you remember me? In memoriam ... the best of the worst Trump pundits https://t.co/J04tJ28yfG
iamtherebel5981|RiotTenMusic|0.6597|0.0|0.722|0.278|RT @RiotTenMusic: 2 things I like more than Trump &amp; Clinton (would probably make better presidents too)  https://t.co/MpfWQ9k4MF
iamtherebel5981|twitter|0.6597|0.0|0.722|0.278|RT @RiotTenMusic: 2 things I like more than Trump &amp; Clinton (would probably make better presidents too)  https://t.co/MpfWQ9k4MF
JTrittini|samkalidi|0.0|0.0|1.0|0.0|RT @samkalidi: @samkalidi Melania Trump be like... https://t.co/8yv9M8ekTA
JTrittini|twitter|0.0|0.0|1.0|0.0|RT @samkalidi: @samkalidi Melania Trump be like... https://t.co/8yv9M8ekTA
CurryForMVP|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
jesseszn_|brooke_hawley5|0.0|0.0|1.0|0.0|RT @brooke_hawley5: Cant wait until Barack Obama is finally out of office tomorrow and Donald Trump is our next precedent #MakeAmericaGrea
SicilianIrish02|Breaking911|-0.6705|0.256|0.744|0.0|RT @Breaking911: PHOTOS: Trump Tower Surrounded By Dump Trucks Filled With Sand To Edge Against Attacks - TMZ https://t.co/DxcqUSuIXT
SicilianIrish02|twitter|-0.6705|0.256|0.744|0.0|RT @Breaking911: PHOTOS: Trump Tower Surrounded By Dump Trucks Filled With Sand To Edge Against Attacks - TMZ https://t.co/DxcqUSuIXT
asahi_azumane|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
asahi_azumane|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
spalienaceship|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Kota_J_S|NathanZed|0.5719|0.0|0.866|0.134|RT @NathanZed: if trump wins im moving to my grandmas house. she still live in america this don't got anything to do with politics I just m
Juanivinazv|ClaireCW76|0.626|0.0|0.687|0.313|RT @ClaireCW76: @DonaldJTrumpJr @realDonaldTrump  WE'RE PRAYING for you President Trump!!! 
jsea226|MagicRoyalty|0.8225|0.0|0.714|0.286|RT @MagicRoyalty: WOW: another proof of #VoterFraud!! Machine refuses to allow vote for Trump!!RT b/c Media will never report this! http
iamronaldpaul|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @Slate @votecastr @LilSteelerGirl @DebAlwaystrump @Kerri1111 TRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLID
BestFrenz|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
BestFrenz|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
onegirlcircus|druchunas|0.7506|0.0|0.73|0.27|"RT @druchunas: Dear Media, after today, please resist the urge to ever publish or produce a story about Donald Trump again. Thank you, Sane"
kitkit22|realDonaldTrump|0.0|0.0|1.0|0.0|@realDonaldTrump TRUMP TRAIN GEORGIA https://t.co/BJ6T4DWe10
kitkit22|twitter|0.0|0.0|1.0|0.0|@realDonaldTrump TRUMP TRAIN GEORGIA https://t.co/BJ6T4DWe10
Mahoney2John|bluehand007|0.0|0.0|1.0|0.0|@bluehand007 president trump
_Nayeelyy|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
_Nayeelyy|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
nemotoad|bigbadjoe21|0.5994|0.122|0.627|0.251|RT @bigbadjoe21: How fitting Trump started his campaign with Latino hate and Latinos can shut him down I love it poetic justice https://t.c
nemotoad||0.5994|0.122|0.627|0.251|RT @bigbadjoe21: How fitting Trump started his campaign with Latino hate and Latinos can shut him down I love it poetic justice https://t.c
slaykingirwin|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
dashiemama|TheRyanParker|0.4019|0.0|0.863|0.137|RT @TheRyanParker: These #TrumpCake memes are going to help us all get through the night: https://t.co/oiuXDIrSf9 #electionday https://t.co
dashiemama|hollywoodreporter|0.4019|0.0|0.863|0.137|RT @TheRyanParker: These #TrumpCake memes are going to help us all get through the night: https://t.co/oiuXDIrSf9 #electionday https://t.co
chrgdup1973|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
Pegasis38|michaeljohns|0.0|0.0|1.0|0.0|RT @michaeljohns: #Pennsylvania:Polls close at 8pm ET (in one hour). Find your polling location here:https://t.co/5wa27WJ8z1#TrumpPA
Pegasis38|pavoterservices|0.0|0.0|1.0|0.0|RT @michaeljohns: #Pennsylvania:Polls close at 8pm ET (in one hour). Find your polling location here:https://t.co/5wa27WJ8z1#TrumpPA
OriginalVader1|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: RCP average in Indiana has Trump up 10.  He is currently up close to 50!!!  Monster vote?  Crossovers?
tennisballbondi|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
tennisballbondi|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
BustosBella|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
LongBlackLine|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
ManikRathee|costareports|0.0|0.0|1.0|0.0|"RT @costareports: On the phone w/ Giuliani. He just left Trump's apt. Said Trump is ""watching everything even tho I'm telling him not to."""
TheUSARocks|mitchellvii|0.2177|0.137|0.684|0.179|RT @mitchellvii: So was Trump winning CO and conveniently every voting machine in the state broke?
alex_saxton21|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
alex_saxton21|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
_3Digital|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_3Digital|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
thetailchaser|MWellerFX|-0.1877|0.088|0.912|0.0|"@MWellerFX @ForexLive @votecastr I saw earlier didnt understand, honestly. But compared to 2012's thresholds, Trump is ahead all but FL"
__shi_ge__|sharonclott|-0.6249|0.231|0.769|0.0|RT @sharonclott: More footage of the topless protest against Trump at my polling station. Two women arrested. #Election2016 https://t.co/bu
__shi_ge__|t|-0.6249|0.231|0.769|0.0|RT @sharonclott: More footage of the topless protest against Trump at my polling station. Two women arrested. #Election2016 https://t.co/bu
FM1888|Bro_Pair|0.0258|0.0|0.936|0.064|@Bro_Pair  I think my ceaseless tweeting about the election to my 140 porn-bot followers has prevented a Trump victory.
Haley_Greentree|rnlisa64|0.0|0.0|1.0|0.0|RT @rnlisa64: Voted Trump!!! #MAGA https://t.co/FTWASnfuRJ
Haley_Greentree|twitter|0.0|0.0|1.0|0.0|RT @rnlisa64: Voted Trump!!! #MAGA https://t.co/FTWASnfuRJ
michaela__16|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
michaela__16|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Coach_DL|MensHumor|0.0|0.0|1.0|0.0|RT @MensHumor: When bae opens up her DMs. https://t.co/Tg1Ovm54cj https://t.co/zwxhkpvCcC
Coach_DL|viralcrunch|0.0|0.0|1.0|0.0|RT @MensHumor: When bae opens up her DMs. https://t.co/Tg1Ovm54cj https://t.co/zwxhkpvCcC
bxnitvvpplebum_|theGrio|-0.1531|0.096|0.904|0.0|RT @theGrio: That awkward moment when you get booed at your own polling place: https://t.co/IOfOYut1ox https://t.co/VBliiVpBCB
bxnitvvpplebum_|thegrio|-0.1531|0.096|0.904|0.0|RT @theGrio: That awkward moment when you get booed at your own polling place: https://t.co/IOfOYut1ox https://t.co/VBliiVpBCB
james_baumann|FastCompany|0.5574|0.0|0.833|0.167|"RT @FastCompany: 16,000 people say they will point and laugh at Trump Tower in NYC tomorrow https://t.co/De92ytpoHC #ElectionDay #Vote2016"
james_baumann|news|0.5574|0.0|0.833|0.167|"RT @FastCompany: 16,000 people say they will point and laugh at Trump Tower in NYC tomorrow https://t.co/De92ytpoHC #ElectionDay #Vote2016"
CaryFrazee|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
sbca80|TheEconomist|-0.7506|0.39|0.61|0.0|RT @TheEconomist: Donald Trump's reckless foreign policy could unleash chaos https://t.co/kJPHr47hHn https://t.co/VhOjRhE6br
sbca80|economist|-0.7506|0.39|0.61|0.0|RT @TheEconomist: Donald Trump's reckless foreign policy could unleash chaos https://t.co/kJPHr47hHn https://t.co/VhOjRhE6br
Amac_16|immigrant4trump|0.7506|0.0|0.766|0.234|"RT @immigrant4trump: If you make this go viral, Trump will win. It's about 2 minutes that makes the choice in this election crystal clear h"
CollinsLowland|NormOrnstein|0.0|0.0|1.0|0.0|RT @NormOrnstein: Maybe he meant both sides of the Trump family https://t.co/gKWBfNmMhY
CollinsLowland|twitter|0.0|0.0|1.0|0.0|RT @NormOrnstein: Maybe he meant both sides of the Trump family https://t.co/gKWBfNmMhY
AnnieBowl|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
haydeemurillo|Fusion|-0.128|0.113|0.795|0.092|"RT @Fusion: ""Since he's gonna lose, I'm going to go dancing.""Latinas share #ElectionNight predictions at the Nevada store Trump tried &amp; f"
stefanivictor1|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
lunaazul70|t|0.0|0.0|1.0|0.0|"https://t.co/64CmtER4LyLive coverage: Election Day 2016 coverage with Katie Couric, Matt Bai"
Marzhattan|JamilahLemieux|-0.2732|0.087|0.87|0.043|"RT @JamilahLemieux: No matter what happens tonight, the fact that Donald Trump has gotten this far is a stain on America that can't be wash"
StamMashiga|themikvahocker|-0.5859|0.375|0.625|0.0|"I think If Trump loses hes gonna have ""CLINTIN""uous tantrums. @themikvahocker"
Jakearias19|Sofy1202|0.5719|0.0|0.748|0.252|RT @Sofy1202: if Trump wins I'll PayPal everyone $1 that RTs this.
suohuu|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
___anet|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
SianJasper|OwensDamien|-0.561|0.256|0.646|0.099|"RT @OwensDamien: Lets hope the closing shot of this terrible movie is Trump all alone in his gold apartment, realising hes forgotten his"
creditclean9|BarbMuenchen|0.4796|0.0|0.865|0.135|RT @BarbMuenchen: URGENT! Calling all #Florida voters and PanHandle of #Florida voters Get out and vote! Trump campaign calling all voters
styleswannabe|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
styleswannabe|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
marianescobar7|jancarlobg|0.0|0.0|1.0|0.0|RT @jancarlobg: F*ck Donald Trump 
waterfunus43|DonaldJTrumpJr|-0.3595|0.098|0.902|0.0|RT @DonaldJTrumpJr: Media elites have done everything they can to stop Trump. WE THE PEOPLE will rise up and take back America! #Trump #Ele
GarrulousGooner|WetherspoonsUK|0.4199|0.0|0.866|0.134|RT @WetherspoonsUK: Choosing between Trump and Clinton for President is like choosing between Wetherspoons and Yates's for your wedding!#E
Meganwiley204|DonaldJTrumpJr|-0.3595|0.098|0.902|0.0|RT @DonaldJTrumpJr: Media elites have done everything they can to stop Trump. WE THE PEOPLE will rise up and take back America! #Trump #Ele
VeilRising13EA|JOMainEvent|0.7456|0.0|0.776|0.224|RT @JOMainEvent: It is the Trump supporters who are the NEW REPUBLICAN PARTY. These landslide victories you see in Senate races is our doin
iamvega1982|ddale8|0.0|0.0|1.0|0.0|"RT @ddale8: Man. Trump, just now, falsely claims that people voting Republican are having their votes switched to Democrats: https://t.co/1"
iamvega1982|twitter|0.0|0.0|1.0|0.0|"RT @ddale8: Man. Trump, just now, falsely claims that people voting Republican are having their votes switched to Democrats: https://t.co/1"
LynnInCA|McDanielJustine|0.0|0.0|1.0|0.0|RT @McDanielJustine: Toomey says he voted for trump
_KrissyGomez|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
CarolBurnett3|twitter|0.7713|0.0|0.599|0.401|"Yes, may we remember who really loves the American People...Trump 2016 https://t.co/dC8sdcNN2K"
jamieross11|jamieross11|-0.8334|0.282|0.718|0.0|"@jamieross11 but while is Clinton is undoubtably corrupt, Trump mighty we'll be the most vile thing on this planet. Tough break 'Murica."
luntaarong|JYSexton|-0.6874|0.294|0.706|0.0|"RT @JYSexton: If Trump freaks out and destroys the Trump Cake, this whole thing still wasn't worth it but..."
swimlife_|jamesmichael|-0.2732|0.084|0.916|0.0|RT @jamesmichael: s/o to this golden moment where Trump let us all know that he doubted his own wife would vote for him. https://t.co/rDdUt
swimlife_|t|-0.2732|0.084|0.916|0.0|RT @jamesmichael: s/o to this golden moment where Trump let us all know that he doubted his own wife would vote for him. https://t.co/rDdUt
iridescentnoir|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
iridescentnoir|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
niahbiah_|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
niahbiah_|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
jskylerinc|HCwrites|-0.5267|0.267|0.631|0.102|RT @HCwrites: A Trump supporter in Florida was just arrested after pulling gun outside polling place https://t.co/dBpQYpPJcb
jskylerinc|usuncut|-0.5267|0.267|0.631|0.102|RT @HCwrites: A Trump supporter in Florida was just arrested after pulling gun outside polling place https://t.co/dBpQYpPJcb
scott006648|WDFx2EU8|-0.4588|0.2|0.8|0.0|RT @WDFx2EU8: Nevada Poll Workers Break Law: Caught Wearing 'Defeat Trump' T-Shirts https://t.co/YaoZoaCPrj
scott006648|thegatewaypundit|-0.4588|0.2|0.8|0.0|RT @WDFx2EU8: Nevada Poll Workers Break Law: Caught Wearing 'Defeat Trump' T-Shirts https://t.co/YaoZoaCPrj
mayadiez|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Purrcival|mjbeckel|-0.4019|0.109|0.891|0.0|"RT @mjbeckel: Who was Trump's biggest ally on the TV airwaves in 2016? The NRA, which aired ~14,000 ads in battleground states https://t.co"
Purrcival|t|-0.4019|0.109|0.891|0.0|"RT @mjbeckel: Who was Trump's biggest ally on the TV airwaves in 2016? The NRA, which aired ~14,000 ads in battleground states https://t.co"
bitchofsaigon|twitter|0.0|0.0|1.0|0.0|I lowkey think she's voting Trump bUTIDK https://t.co/MCbgsx8S7k
DaCrunch|RawStory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
DaCrunch|rawstory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
cisppetta|ReturnofRV|-0.4939|0.132|0.868|0.0|"RT @ReturnofRV: Media will call Florida in order to try to depress Trump turnout in Colorado, Michigan, Nevada. Don't fall for it."
aracelyloll|Ryan23675317|0.4767|0.098|0.675|0.227|RT @Ryan23675317: Just in case trump wins I'm latin btw I'll miss yall
TherealMelHall|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
TherealMelHall|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
sf49ersfan5249|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: #Florida:Trump 48 (+4)Clinton 44Johnson 2#Ohio:Trump 49% (+5)Clinton 44%Johnson 2@trfgrp (R) Poll 10/24-26h
TheMadHessian|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
TheMadHessian|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Solo_Conectate|mashable|0.3612|0.0|0.839|0.161|Trump's website had a glitch that would make it say whatever you'd like https://t.co/zPzH9YbPEH #SoloConectate
teamcombover16|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
3e240ec6b65941b|marshawright|0.0|0.0|1.0|0.0|RT @marshawright: KENTUCKY EARLY RESULTS EXIT POLLSEARLY LEADS POTUS ALERTTRUMP 67.4%CLINTON 28.5%#ElectionNight #electionday #IVOT
annyglop23|Latina_pe|0.0|0.0|1.0|0.0|RT @Latina_pe: Boca de urna- New Hampshire: Donald Trump: 52% Hillary Clinton: 41% #EleccionesEEUU #ElectionDay https://t.co/uhnyqN3ZuC
annyglop23|twitter|0.0|0.0|1.0|0.0|RT @Latina_pe: Boca de urna- New Hampshire: Donald Trump: 52% Hillary Clinton: 41% #EleccionesEEUU #ElectionDay https://t.co/uhnyqN3ZuC
Mvrtial|twitter|0.0|0.0|1.0|0.0|Explain why Clinton &gt; Trump https://t.co/4cxWG5U2dH
Celticlassy10|GissiSim|0.5106|0.0|0.708|0.292|RT @GissiSim: Trump cake memes going strong #ElectionNight https://t.co/oxjcKdQxSl
Celticlassy10|twitter|0.5106|0.0|0.708|0.292|RT @GissiSim: Trump cake memes going strong #ElectionNight https://t.co/oxjcKdQxSl
Cherokee44|thehill|-0.5719|0.258|0.657|0.085|RT @thehill: Trump camp already blaming top Republicans for possible Trump loss before polls close https://t.co/k1feERz6tE https://t.co/qsA
Cherokee44|thehill|-0.5719|0.258|0.657|0.085|RT @thehill: Trump camp already blaming top Republicans for possible Trump loss before polls close https://t.co/k1feERz6tE https://t.co/qsA
john_zealand|Democrat_4Trump|0.0|0.0|1.0|0.0|RT @Democrat_4Trump: &lt;1% votes counted and Trump is leading as per Fox News. If you see #VOTERFRAUD call the POLICE ASAP. Keep watch folks.
MalaineGill|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
MalaineGill|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
HigashiNY|dril|0.0|0.0|1.0|0.0|RT @dril: if you ask me this election could end about 100 different ways:1) trump gets 0% of the vote2) trump gets 1% of the vote3) trum
NorthernTails1|betioserrano|0.2942|0.0|0.856|0.144|RT @betioserrano: Machine Refuses to Allow Vote For Trump in Pennsylvania! #VoterFraud #ElectionDay https://t.co/QPArM5z9bj
NorthernTails1|twitter|0.2942|0.0|0.856|0.144|RT @betioserrano: Machine Refuses to Allow Vote For Trump in Pennsylvania! #VoterFraud #ElectionDay https://t.co/QPArM5z9bj
mcwhirter81|Thomas1774Paine|-0.3612|0.122|0.878|0.0|RT @Thomas1774Paine: #Trump Voters Complain Their Votes Locked Out of Electronic Voting Machines in New York **RT**RT**RT** #voterfraud htt
Delvin_Leon|TheHoodVines|0.8126|0.0|0.575|0.425|RT @TheHoodVines: Me if Trump wins vs. Me if Hilary wins https://t.co/i2n70DTcvi
Delvin_Leon|twitter|0.8126|0.0|0.575|0.425|RT @TheHoodVines: Me if Trump wins vs. Me if Hilary wins https://t.co/i2n70DTcvi
sapersteinjake1|Kylefeldman|0.0|0.0|1.0|0.0|RT @Kylefeldman:  TRUMP TRAIN  https://t.co/xO25CHzq6l
sapersteinjake1|twitter|0.0|0.0|1.0|0.0|RT @Kylefeldman:  TRUMP TRAIN  https://t.co/xO25CHzq6l
CherishedSolace|mmfafa|0.5267|0.103|0.647|0.25|"RT @mmfafa: Fox News just played the ""Blame Russia"" Card...Trump MUST be winning. @mitchellvii @Cernovich @AwesomeIva @StefanMolyneux @Pris"
lildg54|danmericaCNN|0.6037|0.0|0.829|0.171|"RT @danmericaCNN: Khizr Khan to Donald Trump at Clinton's NH event: ""Thankfully, Mr. Trump, this isnt your America."" - Full: https://t.co/"
lildg54|t|0.6037|0.0|0.829|0.171|"RT @danmericaCNN: Khizr Khan to Donald Trump at Clinton's NH event: ""Thankfully, Mr. Trump, this isnt your America."" - Full: https://t.co/"
ButlersEmporium|theguardian|0.0|0.0|1.0|0.0|The Guardian view on Americas choice: Dont vote for Trump. Elect Clinton | Editorial https://t.co/qFbMG3lL0u
berkleyparton|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
smp0711|Gop42016|0.2263|0.095|0.748|0.156|RT @Gop42016: Liberal Bias: Reuters Pulls Polls Showing Huge Trump Surge https://t.co/cGT9cyMFGQ https://t.co/4mhQZbBWVK
smp0711|conservativeread|0.2263|0.095|0.748|0.156|RT @Gop42016: Liberal Bias: Reuters Pulls Polls Showing Huge Trump Surge https://t.co/cGT9cyMFGQ https://t.co/4mhQZbBWVK
hannah_grace_00|jasminewathen19|-0.1531|0.086|0.856|0.059|"RT @jasminewathen19: my 8 year old brother just said ""i want trump to be president because i wanna climb a wall"" im in tears"
BreMichelleee14|HillaryClinton|0.128|0.177|0.622|0.201|"RT @HillaryClinton: Today, let's show the world that love will always trump hate. https://t.co/jfd3CXu1CS https://t.co/a7FXGtAfiG"
BreMichelleee14|hillaryclinton|0.128|0.177|0.622|0.201|"RT @HillaryClinton: Today, let's show the world that love will always trump hate. https://t.co/jfd3CXu1CS https://t.co/a7FXGtAfiG"
OohSterling_|qveen_evelyn|0.3612|0.0|0.873|0.127|RT @qveen_evelyn: If Donald Trump wins.. White people about to think this the 1800's again yeah come side ways if you want to get yo as
scottthong|mitchellvii|0.5719|0.0|0.829|0.171|"RT @mitchellvii: Trump now up 23,000 including Indies in Pinellas County, FL.  In 2012, Obama won this by 26,000."
GreysExorcist|PrimmyRBLX|-0.34|0.338|0.5|0.163|RT @PrimmyRBLX: Pls let trump lose
lewlove123|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
lewlove123|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
anna_rayann|DepressedDarth|0.0|0.0|1.0|0.0|RT @DepressedDarth: Who did you vote for?Retweet for VaderLike for Trump https://t.co/G47xzm8LWV
anna_rayann|twitter|0.0|0.0|1.0|0.0|RT @DepressedDarth: Who did you vote for?Retweet for VaderLike for Trump https://t.co/G47xzm8LWV
808gardeniaG|BarbMuenchen|0.6006|0.0|0.769|0.231|RT @BarbMuenchen: MICHIGAN IS VOTING TRUMP IN HUGE NUMBERS!!  LANDSLIDE VICTORY! https://t.co/QzjPZXtg6H via @wordpressdotcom
808gardeniaG|themarshallreport|0.6006|0.0|0.769|0.231|RT @BarbMuenchen: MICHIGAN IS VOTING TRUMP IN HUGE NUMBERS!!  LANDSLIDE VICTORY! https://t.co/QzjPZXtg6H via @wordpressdotcom
lynn_carleton|pqpolitics|-0.128|0.108|0.803|0.088|RT @pqpolitics: Nato puts 300k troops on 'high alert' as tensions with Russia mount. Which countries would trump let Putin invade? https://
lynn_carleton||-0.128|0.108|0.803|0.088|RT @pqpolitics: Nato puts 300k troops on 'high alert' as tensions with Russia mount. Which countries would trump let Putin invade? https://
PabloPicapiedr7|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
angelrains|video|0.4019|0.0|0.649|0.351|Donald Trump Election Watch Party | https://t.co/xvzumoMGWs
GreyMadison|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
trudybush|AnupKaphle|0.0|0.0|1.0|0.0|RT @AnupKaphle: VIDEO: Donald Trump gets booed as he arrives at his polling place. https://t.co/CJcmBIt9Zl
trudybush|twitter|0.0|0.0|1.0|0.0|RT @AnupKaphle: VIDEO: Donald Trump gets booed as he arrives at his polling place. https://t.co/CJcmBIt9Zl
GAGOPGirl|trfgrp|0.0|0.0|1.0|0.0|"RT @trfgrp: Our projection: Trump 306 Clinton 223 w/CO, VA &amp; WI possibly breaking Trump as ""hidden voter"" #trumptiderolls https://t.co/u34D"
GAGOPGirl|t|0.0|0.0|1.0|0.0|"RT @trfgrp: Our projection: Trump 306 Clinton 223 w/CO, VA &amp; WI possibly breaking Trump as ""hidden voter"" #trumptiderolls https://t.co/u34D"
ItsEcortez|Dianely__alee|0.7351|0.0|0.64|0.36|RT @Dianely__alee: If trump wins I'ma show up to my rancho like https://t.co/RKyulIfdLd
ItsEcortez|twitter|0.7351|0.0|0.64|0.36|RT @Dianely__alee: If trump wins I'ma show up to my rancho like https://t.co/RKyulIfdLd
Kaleymichellea|Buzzthegreatt|0.6249|0.138|0.513|0.349|RT @Buzzthegreatt: I just know Trump gon say something funny when he lose lmao 
juddgreenstein|twitter|0.0|0.0|1.0|0.0|That Trump cake is Batman Walken https://t.co/tS3wdElbat
ChiefMya|haylealsina|-0.8934|0.342|0.588|0.07|@haylealsina shit I'd rather Hillary . Because trump just hell naw . He racist af . Like tf ... And if he become president it's over for us
taaycozart|BOOMINCA|-0.5994|0.206|0.794|0.0|"RT @BOOMINCA: ""*BREAKING NEWS*: Donald Trump and Hilary Clinton both die after their planes collide""America: https://t.co/HjnQMEh6VD"
taaycozart|twitter|-0.5994|0.206|0.794|0.0|"RT @BOOMINCA: ""*BREAKING NEWS*: Donald Trump and Hilary Clinton both die after their planes collide""America: https://t.co/HjnQMEh6VD"
InsaneTrvpper|kiingdarry|0.6249|0.102|0.665|0.232|"RT @kiingdarry: all y'all saying y'all not voting b/c y'all don't believe in Hillary nor Trump, if trump wins Y'ALL BETTER NOT COMPLAIN ABO"
mowser1970|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
fiddyshadz|AndrewKragie|0.3818|0.112|0.683|0.205|"RT @AndrewKragie: Another charmer: man in Kiss outfit, Trump face &amp; hat chants Trump's name as man arrested for sign placement https://t.co"
fiddyshadz|t|0.3818|0.112|0.683|0.205|"RT @AndrewKragie: Another charmer: man in Kiss outfit, Trump face &amp; hat chants Trump's name as man arrested for sign placement https://t.co"
KatieMullock|LeafyIsHere|0.4238|0.139|0.589|0.272|"RT @LeafyIsHere: If Trump wins I'll release nudes, not a joke"
sinncityx|localblactivist|0.0|0.0|1.0|0.0|RT @localblactivist: This correlates to the many instances Trump has pointed out Hillarys war-mongering activities and wall street ties.
mrstiggers1959|RealBenCarson|0.68|0.057|0.697|0.246|@RealBenCarson thank you for all your hard work Mr Carson America willing be rewarded with Mr Trump as our President!
sivanzustin|politico|0.6374|0.0|0.588|0.412|so trump is winning so far??? https://t.co/IoLyxD2sJx
saltprincess77|joelpollak|0.4019|0.0|0.838|0.162|RT @joelpollak: Trump Fans Sing Star-Spangled Banner in Front of Victory Party https://t.co/wVlNFT9hzp via @BreitbartNews
saltprincess77|breitbart|0.4019|0.0|0.838|0.162|RT @joelpollak: Trump Fans Sing Star-Spangled Banner in Front of Victory Party https://t.co/wVlNFT9hzp via @BreitbartNews
kirkbull|dale_bernadette|-0.4574|0.166|0.834|0.0|RT @dale_bernadette: @seanhannity Pennsylvania voters complained of their vote 2 Trump wld switch to Hillary. Frauding again?!
lorna2105|DanielCameron3|0.7184|0.0|0.769|0.231|"RT @DanielCameron3: If Trump wins, when he makes his victory speech I urge @MichelleObama to run behind and scant him. Please retweet. #USE"
KlNDAKELS|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
JordanKingOfOoo|ImDontai|0.0|0.0|1.0|0.0|RT @ImDontai: Told my mom I'm voting for Donald Trump...listen to her reaction  https://t.co/EEa4qQSyKO
JordanKingOfOoo|twitter|0.0|0.0|1.0|0.0|RT @ImDontai: Told my mom I'm voting for Donald Trump...listen to her reaction  https://t.co/EEa4qQSyKO
REAL_Cey_zar|guaptimus_prime|0.0|0.0|1.0|0.0|"RT @guaptimus_prime: There's a ""Trump / Pence"" sign here and this woman in front of me in line TO VOTE just said ""I didn't know Trump's las"
AmBricholas|angryblackhoemo|-0.3595|0.122|0.878|0.0|"RT @angryblackhoemo: white liberals: ""I'm voting for Clinton to stop Trump's racism!""Black people: *lists out ways Hillary's also a racis"
breelieber|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
breelieber|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
nancyl367|Kotcha301|0.4442|0.0|0.867|0.133|RT @Kotcha301: @mitchellvii inside sources are saying Trump landslide. Get out and vote folks. They can't steal this from US!
ELZUNIA79|YoungDems4Trump|0.8126|0.0|0.641|0.359|@YoungDems4Trump @Darren32895836 please vote Trump he is a good man he will take care of us and the country
Highfivemike|USElection_16|-0.4939|0.144|0.856|0.0|Scary to think that a more credible politician could run for president by articulating Trump's policies in four years time @USElection_16
briannag21|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
briannag21|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
electricpac|DiamondandSilk|0.0|0.0|1.0|0.0|"RT @DiamondandSilk: .@realDonaldTrump is Americans only Choice.  Blacks, whites, Hispanics, Asian, Latinos  Vote, Vote, Vote. ......Vote Tr"
imSharna|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
tdotsavage00|twitter|0.8225|0.0|0.591|0.409|When u wanted hillary to win but Trump might actually win #distewmuch #andimeanthat https://t.co/TI9ktXGH4N
starsbombb|3824Miguel|0.0516|0.232|0.526|0.241|"RT @3824Miguel: If Trump wins, i'm playing the longest game of Hide and Seek real shit "
bajanfocus|dib_bee|0.4019|0.0|0.847|0.153|@dib_bee Fact that Trump is a leading candidate of a major US party speak volumes about the country
drunksalamander|brujaaverde|-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
drunksalamander||-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
SaraLindaSimmon|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
ThePJHead|TrumpCardDeck|0.0|0.0|1.0|0.0|RT @TrumpCardDeck: SOURCE: https://t.co/JROXflV0Zy EVIDENCE OF MACHINE MALFUNCTION/FRAUD. Also why is Trump beneath Jill Stein &amp; Gary Johns
ThePJHead|facebook|0.0|0.0|1.0|0.0|RT @TrumpCardDeck: SOURCE: https://t.co/JROXflV0Zy EVIDENCE OF MACHINE MALFUNCTION/FRAUD. Also why is Trump beneath Jill Stein &amp; Gary Johns
Ligi20|CNN|0.25|0.0|0.895|0.105|"RT @CNN: Donald Trump peeked at Melania's ballot, and Twitter had some jokes. Big league. https://t.co/673JwvzlDn #ElectionDay https://t.co"
Ligi20|cnn|0.25|0.0|0.895|0.105|"RT @CNN: Donald Trump peeked at Melania's ballot, and Twitter had some jokes. Big league. https://t.co/673JwvzlDn #ElectionDay https://t.co"
MaureenPeronne|KellyannePolls|0.7096|0.0|0.781|0.219|RT @KellyannePolls: Trump Campaign &amp; RNC @Reince hand in glove. This is about GOP elected officials bragging they voted 3rd party or skippe
NorwayForTrump|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
StLouis_13|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
StLouis_13|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
califsurvivor|Democrat_4Trump|0.0|0.0|1.0|0.0|RT @Democrat_4Trump: &lt;1% votes counted and Trump is leading as per Fox News. If you see #VOTERFRAUD call the POLICE ASAP. Keep watch folks.
enfingercolton2|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: If KY holds anywhere near current levels, Trump will outperform polls there by 35 points."
cesarcarvalho2|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
JankowiakJoAnn|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
whatever_nvm|cihaim|-0.6071|0.386|0.409|0.206|RT @cihaim: GUYS IM CRYING IM SO SCARED THAT TRUMP MIGHT WIN
JohnWalsh001|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
amswank|micahwavee|0.802|0.0|0.647|0.353|RT @micahwavee: I think Hillary &amp; Trump supporters alike can at least agree that Branstad needs to go lol.
cheeseman6697|DonaldJTrumpJr|0.8398|0.0|0.69|0.31|"RT @DonaldJTrumpJr: Please watch and share this. Vote now to take back America! ""Freedom is never more than one generation away from exti"
emmasmommy710|NorahODonnell|0.25|0.0|0.923|0.077|"RT @NorahODonnell: Trump manager @KellyannePolls tells me: ""we are banking on big day of vote in NC, FL, and NV"" to offset Dem EV advantage"
d_edmonds42|jaleighhh_|0.0|0.0|1.0|0.0|RT @jaleighhh_: Trump trump trump
ffforme59|realDonaldTrump|0.3612|0.0|0.848|0.152|RT @realDonaldTrump: 'What I Like About Trump ... and Why You Need to Vote for Him'https://t.co/6rVuDUehZq
itsdjamp|danielgotskillz|0.2732|0.0|0.792|0.208|RT @danielgotskillz: When i see a female Trump supporter lmaoo https://t.co/GjnbUM8Mc2
itsdjamp|twitter|0.2732|0.0|0.792|0.208|RT @danielgotskillz: When i see a female Trump supporter lmaoo https://t.co/GjnbUM8Mc2
northcoastblog|chrislhayes|0.0|0.0|1.0|0.0|"RT @chrislhayes: After waiting until almost *literally* the last moment, Toomey votes and says he voted for Trump."
htall22|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
england_donald|england_donald|0.0|0.0|1.0|0.0|RT @england_donald: A man jumped into action Monday when he spotted a woman grabbing a Donald Trump campaign sign from side of highway. htt
jxkesy|brujaaverde|-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
jxkesy||-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
EnriqueE15|jordanbrak|0.0772|0.0|0.944|0.056|RT @jordanbrak: Donald Trump is a reminder that you should just apply for that job you want even if you don't have experience #ElectionNight
Leeeesliee|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
Leeeesliee|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
thatsk_|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
thatsk_|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
MarkellaUvarova|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
MarkellaUvarova|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
NarryPotter98|drewjustinrauhl|0.0516|0.189|0.566|0.245|RT @drewjustinrauhl: It's idiots like her who support the racist and sexist Donald trump https://t.co/42mlEpShZC
NarryPotter98|twitter|0.0516|0.189|0.566|0.245|RT @drewjustinrauhl: It's idiots like her who support the racist and sexist Donald trump https://t.co/42mlEpShZC
awe_rare|ollaollu|0.0|0.0|1.0|0.0|"RT @ollaollu: Hillary: 67,223 votes (29.1%)Trump: 154,176 votes (66.8%)LIVE 6:57:09 PM ET"
mmrobins|wbruce|0.4753|0.083|0.743|0.174|"@wbruce Hey I think 99 Bananas is delicious with hot chocolate!  My trump cocktail will be 2 parts whiskey, 1 part tears"
Dred1994|moenjonh|0.6835|0.137|0.563|0.3|RT @moenjonh: @NeilTurner_ @cindygarrett14 HEADS UP!!#MSM TO MAKE IT LOOK LIKE TRUMP WINNING - SO WE STOP VOTING!!KEEP VOTING https://t.
Dred1994||0.6835|0.137|0.563|0.3|RT @moenjonh: @NeilTurner_ @cindygarrett14 HEADS UP!!#MSM TO MAKE IT LOOK LIKE TRUMP WINNING - SO WE STOP VOTING!!KEEP VOTING https://t.
Canadian_Shield|Canadian_Shield|0.6124|0.0|0.643|0.357|"@Canadian_Shield: Well, it's official... Trump is President. Thanks, @CNN /s #Election2016"
j_holste|Kaladious|0.0|0.0|1.0|0.0|RT @Kaladious: BREAKING : Only Public Poll that Correctly Called Brexit Predicts Trump Victory https://t.co/lZJRowJIMD
j_holste|truthfeed|0.0|0.0|1.0|0.0|RT @Kaladious: BREAKING : Only Public Poll that Correctly Called Brexit Predicts Trump Victory https://t.co/lZJRowJIMD
babyybry|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
babyybry|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
hertbrknsamurai|MikeGrunwald|-0.6818|0.265|0.64|0.094|"RT @MikeGrunwald: 5. He doesn't like that Trump is crude and a former D. But he'll give Trump a pass. ""A wise man changes his mind. A fool"
Peep_Judy|AdelleNaz|0.0|0.0|1.0|0.0|"RT @AdelleNaz: Star-Spangled Banner being sung by diverse group of Americans in front of #HiltonMidtown, where Trump-Pence ElectionNight pa"
szymborskafiend|samsteinhp|-0.4767|0.129|0.871|0.0|RT @samsteinhp: Trump on Fox News this morning says he will have spent $100 million in total. Wrong till the last day
Citizen4NYC|nytimes|-0.4215|0.141|0.859|0.0|"@nytimes Bush v Gore was December 12.  This will be same unless Trump crushed in Fl, OH, &amp; PA."
a_mamii6|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
LindaLouJones13|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
scr385w|NRO|0.0|0.0|1.0|0.0|"RT @NRO: Early Exit Polls: Trump Opens YUGE Gap between College-Educated, Non-College-Educated Whiteshttps://t.co/ADpCNhYfiC #ElectionNight"
daout1aw|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
drafthorse2012|mitchellvii|0.34|0.0|0.893|0.107|"RT @mitchellvii: I expect Trump to win KY and IN, but not by 50 points.  We'll see if anything near that holds."
Shade58b|mitchellvii|0.7998|0.0|0.736|0.264|RT @mitchellvii: The last RCP Poll had Trump winning KY by 17.  He is currently winning by 52 points.Monster vote?  Dem crossovers?
linds_|kurteichenwald|0.3612|0.0|0.898|0.102|RT @kurteichenwald: 40. Trump claimed to own 50% of a project when he owned 30%. His explanation under oath: I always felt like I owned 50
TheValuesVoter|ananavarro|-0.2732|0.087|0.913|0.0|"RT @ananavarro: Hey Nevadans, u know why Trump is suing? To keep Hispanics from polls b/c he knows we're voting against him. Redouble your"
feltinos|ogmaxb|0.25|0.083|0.797|0.12|RT @ogmaxb: Donald Trump saw a boy who was lost in New York and didn't tell anyone.Is this a man we can trust as President? https://t.co/X
feltinos|linkedin|0.25|0.083|0.797|0.12|RT @ogmaxb: Donald Trump saw a boy who was lost in New York and didn't tell anyone.Is this a man we can trust as President? https://t.co/X
abermans|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
MissLiberty1776|DonaldJTrumpJr|0.7644|0.0|0.752|0.248|RT @DonaldJTrumpJr: Young people across the country are rising up voting for Trump. Young democrats have been amazing! Thank you for your v
DavidDarr2|JohnKStahlUSA|-0.8519|0.368|0.632|0.0|RT @JohnKStahlUSA: Undocumented relative charged with killing 10-year-old girl. Still think Trump was wrong? #tcot #ccot #gop #maga  https:
jill19677|coton_luver|-0.0258|0.128|0.749|0.123|RT @coton_luver: A deplorable Trump Fan Just Pulled A Gun On A Black Voter At #Florida Polling Station - https://t.co/EepIioqOJd
jill19677|occupydemocrats|-0.0258|0.128|0.749|0.123|RT @coton_luver: A deplorable Trump Fan Just Pulled A Gun On A Black Voter At #Florida Polling Station - https://t.co/EepIioqOJd
Fomexis|stats_canada|0.4588|0.0|0.824|0.176|RT @stats_canada: Canada is preparing to welcome 150 million American refugees if Trump becomes president
SpencerPolap|FoxNews|0.9296|0.0|0.52|0.48|"@FoxNews Canada needs Trump as well!!! When America is strong, Canada is strong!!! Keep it up Fox News! God Bless America!"
juanzavala67|LouieVRee|-0.8271|0.3|0.636|0.064|RT @LouieVRee: Trump gay as hell if he trying to get rid of all the fine big booty Latina bitches too
killerrays|nathanTbernard|0.1904|0.177|0.602|0.222|"RT @nathanTbernard: @realDonaldTrump Trump will be finished, woo! NO MORE TRUMP! https://t.co/3kkTcBErus"
killerrays|hillaryclinton|0.1904|0.177|0.602|0.222|"RT @nathanTbernard: @realDonaldTrump Trump will be finished, woo! NO MORE TRUMP! https://t.co/3kkTcBErus"
Jayis4_Jasmen|Jayis4_Jasmen|-0.2298|0.241|0.55|0.209|@Jayis4_Jasmen so damn entitled to your own opinions until Trump wins and these racist mfs start rioting in the streets.....
leejooheonanti|naktaofficiaI|0.0516|0.217|0.559|0.224|"RT @naktaofficiaI: donald trump is winning, i thought half of the population in the usa was intelligent and i was wrong, sad"
veroarreguin|latimes|0.0|0.0|1.0|0.0|"The power of an education: To Donald Trump, from the undocumented immigrant who graduated alongside your daughter https://t.co/0QG3KVsBlU"
MeghansMusings|slate|-0.4019|0.153|0.847|0.0|Things Trump could have done instead of wasting his time running for president: https://t.co/04Mst1lAxE via @slate
MeghansMusings|slate|-0.4019|0.153|0.847|0.0|Things Trump could have done instead of wasting his time running for president: https://t.co/04Mst1lAxE via @slate
perkoflaura|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
perkoflaura|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
cutelilbish|twitter|-0.7964|0.333|0.55|0.116|omg read wtf i sed if trump win the earth gonna end cause he gonna fuck sum shit up i voted for #HillaryClinton https://t.co/1Deq5bdRMW
ElectionNewsHQ|twitter|0.0|0.0|1.0|0.0|FOX News Exit Poll among Hispanic Voters:2016Clinton 65%Trump 27%2012Obama 71%Romney 27%#ElectionNight https://t.co/h7BMqULHnD
AvrgeBerenstain|cosmo_8a|0.0258|0.148|0.7|0.152|RT @cosmo_8a: If trump wins and anybody starts a riot let me know I'm trying to get a tv or something
Koipan23|JordanRae_24|0.0|0.0|1.0|0.0|RT @JordanRae_24: a lot of people are tryna vote for trump but the computers are changin it to Hillary 
AdedigbaAdeniy1|washingtonpost|0.3612|0.0|0.839|0.161|"RT @washingtonpost: A Trump presidency would be like Stevie Wonder driving, Stevie Wonder says https://t.co/tLNfxuxYPc"
AdedigbaAdeniy1|washingtonpost|0.3612|0.0|0.839|0.161|"RT @washingtonpost: A Trump presidency would be like Stevie Wonder driving, Stevie Wonder says https://t.co/tLNfxuxYPc"
barbandaaron|twitter|0.4215|0.0|0.851|0.149|"Bring back our rights, jobs, business, amendments, safety, our Healthcare  that is slowly being taken away.America https://t.co/5QE4yy4TAD"
eschwent|carlajo1947|0.0|0.0|1.0|0.0|RT @carlajo1947: REPORTS ARE COMING OUT THAT MICHIGAN VOTING IS CURRENTLY A LANDSLIDE VICTORY FOR TRUMP! https://t.co/eFiVAidr9l
eschwent|twitter|0.0|0.0|1.0|0.0|RT @carlajo1947: REPORTS ARE COMING OUT THAT MICHIGAN VOTING IS CURRENTLY A LANDSLIDE VICTORY FOR TRUMP! https://t.co/eFiVAidr9l
imogen19091|KGBVeteran|0.0|0.0|1.0|0.0|RT @KGBVeteran: Black man flashes Trump #MAGA hat at camera. This is in Cleveland. #ElectionDay https://t.co/qw0NzwHksv
imogen19091|twitter|0.0|0.0|1.0|0.0|RT @KGBVeteran: Black man flashes Trump #MAGA hat at camera. This is in Cleveland. #ElectionDay https://t.co/qw0NzwHksv
lookitslyndseyy|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
betsy1217|RaymondArroyo|-0.3818|0.126|0.874|0.0|RT @RaymondArroyo: The scene outside Trump Tower. Lots of NYPD and dump trucks up and down 5th Ave. https://t.co/wMRy0nHwuC
betsy1217|twitter|-0.3818|0.126|0.874|0.0|RT @RaymondArroyo: The scene outside Trump Tower. Lots of NYPD and dump trucks up and down 5th Ave. https://t.co/wMRy0nHwuC
yugijo|twitter|0.6588|0.0|0.732|0.268|"From the great state of PA, this latina voted for #Trump ! #MAGA https://t.co/1wPZSi4Wpk"
GavinCurnow|KQAnderson|-0.7959|0.336|0.664|0.0|@KQAnderson Holy shit! I just took a pic of some dejected Trump campaigners in the Biloxi McDonalds earlier...
rmontgomery29|worldnetdaily|-0.4588|0.176|0.824|0.0|RT @worldnetdaily: Trump to Savage: 'I used to think real estate was vicious'https://t.co/eEAOnnkYHX@ASavageNation @realDonaldTrump #MAGA
rlpeace|BrockVergakis|-0.2263|0.079|0.921|0.0|RT @BrockVergakis: This Navy veteran took a bus and walked 3 blocks on crutches to vote for Clinton in Norfolk. Says Trump doesn't know mor
VictoriaJoyeuse|RichardBSpencer|0.0|0.0|1.0|0.0|@RichardBSpencer  Most of the rank and file Republicans I have met volunteering are on board with Trump and gradually also with nationalism.
GillandBrad|twitter|0.0|0.0|1.0|0.0|"Trump go California, California go red! https://t.co/m5CmrhKHI1"
creminsmom|JOHNSONSFOOL|-0.4003|0.119|0.881|0.0|@JOHNSONSFOOL If Hillary worked for a bank (any US Company) &amp;  released Confidential Info.... She is fired.... Fire Hillary .... Vote Trump!
twooor|mlissa1|-0.2263|0.142|0.751|0.107|RT @mlissa1: I am a Mexican American that lives in South Texas. Unlike Ana Navarro I clearly heard when Trump said Illegal immigrants. I vo
diabadassss|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
kasstanb|GaryLineker|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
kasstanb|twitter|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
Educate4ward|JasonFebery|0.743|0.109|0.561|0.33|"RT @JasonFebery: Lifelong Republican Ana Navarro: ""It would be sweet, sweet justice if the Hispanic vote defeated Trump tonight."" #Election"
_Zakkery_|FreeMemesKids|-0.1695|0.196|0.804|0.0|"RT @FreeMemesKids: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
stumpyyyyyyy|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Lovely__Souls|caramelthot|-0.1655|0.064|0.936|0.0|"RT @caramelthot: my neighbor just told me someone stole her trump sign last night &amp; i acted all shocked, but little does she know i was the"
jtelofski|shelbyfero|0.6249|0.0|0.769|0.231|RT @shelbyfero: Lol Trump isn't checking that Melania voted for him he's making sure he's doing his ballot right.
RaniaMounir|USATODAY|-0.34|0.13|0.87|0.0|RT @USATODAY: Internet goes crazy over photo of Trump appearing to look at Melania's ballot https://t.co/tmtQvFaeSJ https://t.co/BtkAIIDJFK
RaniaMounir|usatoday|-0.34|0.13|0.87|0.0|RT @USATODAY: Internet goes crazy over photo of Trump appearing to look at Melania's ballot https://t.co/tmtQvFaeSJ https://t.co/BtkAIIDJFK
reinadelreys|rainymondays|0.0|0.0|1.0|0.0|RT @rainymondays: me to 'gays for trump' when i get sent to concentration camps &amp; see them there https://t.co/EI2nKmmPse
reinadelreys|twitter|0.0|0.0|1.0|0.0|RT @rainymondays: me to 'gays for trump' when i get sent to concentration camps &amp; see them there https://t.co/EI2nKmmPse
travestynv|jasonvolack|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
travestynv|twitter|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
vivianbrown21|AsapBasile98|0.0|0.0|1.0|0.0|"RT @AsapBasile98: Today, On #ElectionDay , I voted for : #Trump #HillaryClinton #TrumpPence16 #Election2016 #ClintonVsTrump #electionpoll"
N1GHTR1DE|x0crys|-0.4404|0.195|0.805|0.0|RT @x0crys: if you voted for trump block me and take it personal
shakeiyah_|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
shakeiyah_|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
BJA1021|hrtablaze|0.5399|0.0|0.868|0.132|RT @hrtablaze: CNN reporting that there is record breaking turnout! That is good news for the Trump Train ! First Exit Poll comes out short
ideavator|FreddieCampion|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
ideavator|twitter|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
EmehDR|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
EmehDR|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
r_saunds_21|Philatticus|-0.5719|0.15|0.85|0.0|@Philatticus @SmartySampson too much hate for trump for people to change their minds that happened too late in my opinion possible though
cal_cach3|Pamela_Moore13|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: ENDLESS #VOTERFRAUD!Votes flipped from Trump to Clinton in Pennsylvania. https://t.co/TeDuk0Iu3D
cal_cach3|twitter|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: ENDLESS #VOTERFRAUD!Votes flipped from Trump to Clinton in Pennsylvania. https://t.co/TeDuk0Iu3D
Largr16|darylpfosterpvv|0.0|0.0|1.0|0.0|RT @darylpfosterpvv: Wooow this is Yuuuge!!! Staat Kentucky is poll binnen!! #Trump #CNN https://t.co/za2D656ut9
Largr16|twitter|0.0|0.0|1.0|0.0|RT @darylpfosterpvv: Wooow this is Yuuuge!!! Staat Kentucky is poll binnen!! #Trump #CNN https://t.co/za2D656ut9
SueCFlorida|FredZeppelin12|0.25|0.0|0.895|0.105|RT @FredZeppelin12: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERS. Advantage #Trump. Evening voters are evening voters because t
_tierrrraaaa|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_tierrrraaaa|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
jadejesleighpez|nipplynjh|0.5499|0.094|0.736|0.169|"RT @nipplynjh: No vote = a vote for trump. No one is happy about the options, but you have to do what you have to do to ensure that its any"
Cutellic|maoridays|0.6757|0.0|0.799|0.201|RT @maoridays: if you support trump break the mutual i don't give a fuck how long we've been mutuals break it right now bc i suddenly don't
d6sty|PzFee|0.4404|0.0|0.873|0.127|RT @PzFee: BREAKING NEWS -- Spongebob shot at Trump rally. He was supporting Hillary Clinton and got shot by Plankton. https://t.co/mU8MRF2
d6sty|t|0.4404|0.0|0.873|0.127|RT @PzFee: BREAKING NEWS -- Spongebob shot at Trump rally. He was supporting Hillary Clinton and got shot by Plankton. https://t.co/mU8MRF2
lilwha13|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
lilwha13|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
scummartist|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
scummartist|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
Giography_|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Giography_|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
ay_jay42|TheHoodVines|0.8126|0.0|0.575|0.425|RT @TheHoodVines: Me if Trump wins vs. Me if Hilary wins https://t.co/i2n70DTcvi
ay_jay42|twitter|0.8126|0.0|0.575|0.425|RT @TheHoodVines: Me if Trump wins vs. Me if Hilary wins https://t.co/i2n70DTcvi
O_dealia|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
O_dealia|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
LovinnThaCrew|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
LovinnThaCrew|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
Dj2016djt|debsellsslc|0.5719|0.144|0.608|0.247|RT @debsellsslc: Never Forget those who Risked All 4 our FeedomGod Bless #America #Trump the only Patriot running Loves USA https://
Dj2016djt||0.5719|0.144|0.608|0.247|RT @debsellsslc: Never Forget those who Risked All 4 our FeedomGod Bless #America #Trump the only Patriot running Loves USA https://
mattm4000|juliet0497|0.0|0.0|1.0|0.0|"@juliet0497 ""I Never ran for President.""--Donald Trump 11/9/16."
risejaeb|yugbma|-0.1833|0.24|0.588|0.172|RT @yugbma: im deadass scared like... i do not want to be stuck with trump... god please be with us https://t.co/TqTQvSBirc
risejaeb|twitter|-0.1833|0.24|0.588|0.172|RT @yugbma: im deadass scared like... i do not want to be stuck with trump... god please be with us https://t.co/TqTQvSBirc
leojnalsik|alaskantexanQCT|0.0|0.0|1.0|0.0|RT @alaskantexanQCT: Yo fam heading to Philly with some homies and 2 vans. Gonna take Black Trump voters 2 the polls ALL DAY tomorrow! #MAG
KingKinthehouse|TeenVogue|-0.3595|0.333|0.667|0.0|"RT @TeenVogue: No peeking, Donald! https://t.co/Q2GflxtECB"
KingKinthehouse|teenvogue|-0.3595|0.333|0.667|0.0|"RT @TeenVogue: No peeking, Donald! https://t.co/Q2GflxtECB"
thejenn999|jason_howerton|0.0|0.0|1.0|0.0|RT @jason_howerton: Trump leads Clinton 70.5% to 25.8% in Indiana -- and 68% to 28% in Kentucky with just 2% of the vote in. #ElectionNight
chulabeIIe|Flamemmakins|0.4404|0.0|0.873|0.127|RT @Flamemmakins: @chulabeIIe If I were in Greeley right now I would deadass be driving around town to see these true-life Trump supporters
chrissyrules66|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
pacmann007|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
pacmann007|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
GGIRLYYY_|sogates_|-0.4717|0.305|0.695|0.0|RT @sogates_: if Trump doesn't win president   https://t.co/7tdoCQXHJT
GGIRLYYY_|twitter|-0.4717|0.305|0.695|0.0|RT @sogates_: if Trump doesn't win president   https://t.co/7tdoCQXHJT
He_is_er_man|huntigula|0.4588|0.0|0.846|0.154|RT @huntigula: why do I get the feeling Trump is doing 'the tuck' under that robe like buffalo bill from Silence of the Lambs https://t.co/
He_is_er_man|t|0.4588|0.0|0.846|0.154|RT @huntigula: why do I get the feeling Trump is doing 'the tuck' under that robe like buffalo bill from Silence of the Lambs https://t.co/
_HippieMatthews|divineeCaroline|0.7236|0.0|0.718|0.282|RT @divineeCaroline: You want equality??But you support Trump who wants to deport immigrants who come here searching for equality and freed
miyuwi|CNN|0.0|0.0|1.0|0.0|RT @CNN: This is how close Clinton and Trump will be to each other in Manhattan tonight https://t.co/YPAfWQsye5 #ElectionDay https://t.co/4
miyuwi|cnn|0.0|0.0|1.0|0.0|RT @CNN: This is how close Clinton and Trump will be to each other in Manhattan tonight https://t.co/YPAfWQsye5 #ElectionDay https://t.co/4
lopezzjenn|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
slmorris555|dymaund|-0.5423|0.179|0.821|0.0|"RT @dymaund: at the end of the day, Donald Trump is just a Tv personality with a bad tan....#ImWithHer "
DunkirkDavid|jakerock88|0.7003|0.0|0.746|0.254|@jakerock88 good evening Jake thanks for the follow we need Donald Trump as our president never Hillary @TeamTrump #Election2016
JOETWIT5ST|VincentLombar13|0.0|0.0|1.0|0.0|"RT @VincentLombar13: TRUMP LANDSLIDE      2016""Either we have a country or we don't.""~Donald J Trump https://t.co/IKfvkynfND"
JOETWIT5ST|twitter|0.0|0.0|1.0|0.0|"RT @VincentLombar13: TRUMP LANDSLIDE      2016""Either we have a country or we don't.""~Donald J Trump https://t.co/IKfvkynfND"
Zippittt|mtracey|0.0|0.0|1.0|0.0|"RT @mtracey: Former Sanders delegate from PA sends over this photo: voted Trump, then Democrats down ballot https://t.co/qfwbyhwIFx"
Zippittt|twitter|0.0|0.0|1.0|0.0|"RT @mtracey: Former Sanders delegate from PA sends over this photo: voted Trump, then Democrats down ballot https://t.co/qfwbyhwIFx"
amukamusic|facebook|-0.2228|0.157|0.66|0.183|If you want to know the most racist places in AMERICA...look where Trump is winning! I went to Lapeer MI today... https://t.co/ROywVviabx
TuNaLdO|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
TuNaLdO|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
MackenzieEaton|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
MackenzieEaton|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
wisey_9|Cain_Unable|0.0|0.0|1.0|0.0|"RT @Cain_Unable: I just tried to Vote Trump &amp; the staff wouldn't let me just because I'm ""in Kent"" &amp; ""this is a Tesco self service checkout"
JIndeliclae|brainpicker|-0.6597|0.24|0.702|0.058|"RT @brainpicker: ""Im horrified to watch the bizarre pageant of my nation pretending these two contenders are equivalent."" THIS https://t.c"
JIndeliclae||-0.6597|0.24|0.702|0.058|"RT @brainpicker: ""Im horrified to watch the bizarre pageant of my nation pretending these two contenders are equivalent."" THIS https://t.c"
patrioticwoman3|Trump2016News|0.0|0.0|1.0|0.0|"RT @Trump2016News: Republicans: I know you're all busy WORKING, but don't put off voting at 5PM! Trump never gave up on you; don't give up"
firefly00001101|JohnKStahlUSA|-0.8519|0.368|0.632|0.0|RT @JohnKStahlUSA: Undocumented relative charged with killing 10-year-old girl. Still think Trump was wrong? #tcot #ccot #gop #maga  https:
Dowling_Sam|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
tweIvethirty|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
tweIvethirty|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
luh_lex|Damnimcold32|0.5145|0.088|0.706|0.206|RT @Damnimcold32: If Donald Trump become president nobody better not say shit to me the whole ride back to Mexico or we fighting
caleb_330|Avstvn|-0.1695|0.196|0.804|0.0|"RT @Avstvn: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
Glennard|alliepape|-0.5126|0.182|0.736|0.082|RT @alliepape: A customs official's abuse of power didn't stop this Mission store owner from getting her Trump piatas. https://t.co/vEUQUU
Glennard|t|-0.5126|0.182|0.736|0.082|RT @alliepape: A customs official's abuse of power didn't stop this Mission store owner from getting her Trump piatas. https://t.co/vEUQUU
Nick_Rallis|FauxPelini|-0.5319|0.153|0.847|0.0|RT @FauxPelini: .@realDonaldTrump When I pressed Trump the touchscreen burned my finger and said ERROR &amp; when I pressed Clinton a lady gave
yannlgrnd|riskmaplive|-0.765|0.306|0.694|0.0|RT @riskmaplive: Reports Of Massive Voter Fraud Flood In - Discrimination &amp; Intimidation Aginast Trump Voters https://t.co/EiGwyuuFYj https
yannlgrnd|riskmap|-0.765|0.306|0.694|0.0|RT @riskmaplive: Reports Of Massive Voter Fraud Flood In - Discrimination &amp; Intimidation Aginast Trump Voters https://t.co/EiGwyuuFYj https
buzz|hunterw|0.6249|0.0|0.812|0.188|"RT @hunterw: Media at the Trump party are being kept away from guests in a small area that security described to me as a ""press buffer."""
BryanCusick|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
BryanCusick|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
TheMinerK|TheFunnyVine|-0.0191|0.097|0.903|0.0|RT @TheFunnyVine: Trump and Hillary will never reach this level  https://t.co/9jl1rDKqj7
TheMinerK|vine|-0.0191|0.097|0.903|0.0|RT @TheFunnyVine: Trump and Hillary will never reach this level  https://t.co/9jl1rDKqj7
valeriem03|brujaaverde|-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
valeriem03||-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
Tinasvue|bigboater88|0.4374|0.0|0.879|0.121|RT @bigboater88: Fellow Floridians =  Please don't do anything after work except VOTE TRUMP! Get to your local Poll and VOTE TRUMP! #DrainT
craigmack79|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
craigmack79|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
emileemaeeeh|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
mlynne3|Miami4Trump|0.7003|0.0|0.766|0.234|RT @Miami4Trump: Trump Cares About Inner Cities And Improving Education. He's discussed This For Over 30 YEARS #VoteTrump He Will #MAGA#El
overthetopdani|jamescharles|0.4404|0.0|0.775|0.225|RT @jamescharles: good morning everyone except those voting for Donald Trump
CeletaQ|mms5048|0.0|0.0|1.0|0.0|RT @mms5048: McCain refuses to say he voted for Trump | TheHill - https://t.co/prl08KHWsR
CeletaQ|thehill|0.0|0.0|1.0|0.0|RT @mms5048: McCain refuses to say he voted for Trump | TheHill - https://t.co/prl08KHWsR
sg_scarr|GinaGrif823|0.5904|0.0|0.723|0.277|RT @GinaGrif823: @JOMainEvent @immigrant4trump @CBSNews AND THAT MY FRIENDS IS TRUMP#MAGA
httpmekah|CGGuy44|0.8748|0.0|0.546|0.454|RT @CGGuy44: Good morning! I hope everyone has a blessed day except the 'gays for trump'. https://t.co/xA8zPNnWqw
httpmekah|twitter|0.8748|0.0|0.546|0.454|RT @CGGuy44: Good morning! I hope everyone has a blessed day except the 'gays for trump'. https://t.co/xA8zPNnWqw
patchrhythm|DonnajeanGray3|0.6625|0.0|0.613|0.387|RT @DonnajeanGray3: TRUMP IS WINNING NOW!###LOVE YOU DONALD
Isdat_Morpheus|Scout_Finch|0.0258|0.156|0.684|0.16|RT @Scout_Finch: I will remember you. Will you remember me? In memoriam ... the best of the worst Trump pundits https://t.co/J04tJ28yfG
Isdat_Morpheus|twitter|0.0258|0.156|0.684|0.16|RT @Scout_Finch: I will remember you. Will you remember me? In memoriam ... the best of the worst Trump pundits https://t.co/J04tJ28yfG
willOBell|AmiriKing|0.0|0.0|1.0|0.0|RT @AmiriKing: Idea:Split the U.S. in half.Dems get one side.Reps get one side.Hillary runs your lives.Trump leads ours.#Clinto
bolajoselopez|JordanHyland21|0.3182|0.103|0.7|0.198|RT @JordanHyland21: If Donald Trump wins the election I will Paypal $100 to one person who retweets this. No backing out.
TheUndine3|damaninthearena|0.0|0.0|1.0|0.0|RT @damaninthearena: @Vendetta92429 @antimarxis_ this map is BS!! I'm in southern Cali and in a line of 50+ people; Black White Hispanic As
neurotichealy|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
neurotichealy|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
AguiRuben|SoaRPraizist|0.5719|0.0|0.802|0.198|"RT @SoaRPraizist: If Trump wins the election, I will make artwork for everyone that RTs this tweet"
ryncarnate|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
treyton_davila|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
CharliseAnne|ClarenceJWhite|0.0|0.069|0.863|0.069|RT @ClarenceJWhite: I feel like Trump &amp; Hillary are two divorced parents fighting over custody of us but we kinda just wanna go live with g
Jojo_Lovejoy|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
Jojo_Lovejoy|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
Mafamal|twitter|0.5719|0.0|0.448|0.552|If Trump wins https://t.co/3jwMRvrbzs
GreenBiotechie|chrislhayes|-0.5256|0.159|0.841|0.0|RT @chrislhayes: Trump is already laying the groundwork to contest the legitimacy of the election and it's incredibly dangerous.
carrrrrrina|HillaryClinton|0.128|0.177|0.622|0.201|"RT @HillaryClinton: Today, let's show the world that love will always trump hate. https://t.co/jfd3CXu1CS https://t.co/a7FXGtAfiG"
carrrrrrina|hillaryclinton|0.128|0.177|0.622|0.201|"RT @HillaryClinton: Today, let's show the world that love will always trump hate. https://t.co/jfd3CXu1CS https://t.co/a7FXGtAfiG"
ChristineIs43|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
ayy_its_jaydenn|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
ayy_its_jaydenn|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Nikki_Bitchhh|ShineVista|0.3616|0.148|0.608|0.243|"RT @ShineVista: Prediction: Hillary Clinton wins election, Donald Trump doesn't concede. America riots, &amp; people die. Market crashes. Haram"
Saritrovick|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
Saritrovick|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
NormandinRob|LindaSuhler|0.6776|0.0|0.798|0.202|"RT @LindaSuhler: Your SINGLE VOTE could be the difference between Donald J. Trump winning or not.Whatever it takes, VOTE!!!!#VoteTrump"
njhnetflix|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
nellaenimsaj|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
nellaenimsaj|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
fredgthegreat|GovMikeHuckabee|-0.0516|0.059|0.941|0.0|"RT @GovMikeHuckabee: I personally know both candidates;Have for years; Not hard choice. Neither are perfect-nor am I, but voted Trump w/o h"
NeilShelley|jeremyscahill|0.7269|0.0|0.775|0.225|RT @jeremyscahill: Trump insiders tell me he plans to use shredded copies of his tax returns as confetti tonight after his huge win.
Turboturbulence|KnowbodysTweets|0.2023|0.176|0.621|0.203|RT @KnowbodysTweets: Nah. Now they believe that Trump is the only racist and that the beautiful and fair voting system will eliminate him h
scottthong|mitchellvii|0.7998|0.0|0.736|0.264|RT @mitchellvii: The last RCP Poll had Trump winning KY by 17.  He is currently winning by 52 points.Monster vote?  Dem crossovers?
jeanigum|runningforpizza|0.0|0.0|1.0|0.0|RT @runningforpizza: Hannity is reporting that Florida panhandle residents need to show up for Trump!!!!! Get out and vote!!!! https://t.co
jeanigum|t|0.0|0.0|1.0|0.0|RT @runningforpizza: Hannity is reporting that Florida panhandle residents need to show up for Trump!!!!! Get out and vote!!!! https://t.co
jackelpdubz|Reevellp|0.4019|0.0|0.881|0.119|RT @Reevellp: In #Moscow there is a Trump party in-full swing- pro-Kremlin activists gathered in a bar for the results. Giant portrait of T
waithash|FrankLuntz|-0.1027|0.055|0.945|0.0|RT @FrankLuntz: The turnout in Democratic Philadelphia is so high that it's hard to see Trump overcoming it in the rest of the state.  #Ele
DraftRomney|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: Report: President George W. Bush didn't vote for either Trump, Clinton. #ElectionNight #FoxNews2016 https://t.co/wKkrha8Bqn"
DraftRomney|twitter|0.0|0.0|1.0|0.0|"RT @FoxNews: Report: President George W. Bush didn't vote for either Trump, Clinton. #ElectionNight #FoxNews2016 https://t.co/wKkrha8Bqn"
Vito57817838|Democrat_4Trump|0.0|0.0|1.0|0.0|RT @Democrat_4Trump: Reports are coming out that Michigan voting is currently a landslide victory for Trump. https://t.co/hNgj5Q344w
Vito57817838|twitter|0.0|0.0|1.0|0.0|RT @Democrat_4Trump: Reports are coming out that Michigan voting is currently a landslide victory for Trump. https://t.co/hNgj5Q344w
edenrathore|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
edenrathore|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
stanoliver|LOLGOP|0.0516|0.138|0.714|0.148|RT @LOLGOP: EXIT POLL: 3 in 10 Trump supporters had trouble finding the exit to the polls.
GiselaMDiaz|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
GiselaMDiaz|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
Nexykat|AnonD4ms3l|0.6486|0.057|0.741|0.202|"RT @AnonD4ms3l: Seriously, if you people elect #Pence handpicked errand boy in #Indiana for Gov, or if Trump wins the WH, ima pray for @smo"
allboutendz|GovMikeHuckabee|-0.0516|0.059|0.941|0.0|"RT @GovMikeHuckabee: I personally know both candidates;Have for years; Not hard choice. Neither are perfect-nor am I, but voted Trump w/o h"
comiateerepetia|twitter|0.0|0.0|1.0|0.0|EVERYBODY TRUMP TRUMP TRUMP https://t.co/x0omTPxrZ4
ninability|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
CADOF1|americannewsx|0.4927|0.0|0.862|0.138|"The Trump Trolls are not known for being very bright. Today when they went to vote they learned a new word,... https://t.co/hF146Pa2sl"
TeresaE17|hrtablaze|0.9207|0.0|0.645|0.355|RT @hrtablaze: My Bernie Sanders loving nephew who has been messing with me all election just told me he voted TRUMP !!! WOOT WOOT ! #elect
bigbrownbat|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
bigbrownbat|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
rabbitoh_von|farrm51|-0.3818|0.098|0.902|0.0|RT @farrm51: Karl Rove points out Trump said GWBush knew about &amp; allowed 9/11; lied re WMD; called for impeachment. &amp; wonders why Bush's di
solozaiin|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
solozaiin|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
KevsterYT96|ajbvnks|0.7579|0.0|0.615|0.385|RT @ajbvnks: If you support Donald trump please like this tweet so I can unfollow you
mbaangluuc|DonaldJTrumpJr|0.6114|0.0|0.8|0.2|RT @DonaldJTrumpJr: The fate of America could be determined in the next couple hours. Please do your part. Vote Trump! #MAGA #Election2016
hauserlisa1|bigbare44|0.0|0.0|1.0|0.0|RT @bigbare44: https://t.co/oe3Q6ov9dNTRUMP. TRUMP. TRUMP.
hauserlisa1|t|0.0|0.0|1.0|0.0|RT @bigbare44: https://t.co/oe3Q6ov9dNTRUMP. TRUMP. TRUMP.
VGVG0|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
VGVG0|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
ves_secret|FunnyPicsDepot|0.3612|0.082|0.781|0.138|RT @FunnyPicsDepot: Stop saying if trump wins yall moving out of the country. Stfu yall cant even move outta ya mommas house https://t
ves_secret||0.3612|0.082|0.781|0.138|RT @FunnyPicsDepot: Stop saying if trump wins yall moving out of the country. Stfu yall cant even move outta ya mommas house https://t
brendangill5|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
allencountytp|facebook|0.5719|0.0|0.778|0.222|Based on the Early Vote. Donald Trump has won the state of Indiana. https://t.co/5yCze92gPs
titttaaahh|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
titttaaahh|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
debbiedo58|megynkelly|0.3612|0.0|0.898|0.102|"RT @megynkelly: .@IngrahamAngle: If were going to see a real move for #Trump, its going to have to exist in a state like #Michigan. #El"
_Fer_Ochoa_|jancarlobg|0.0|0.0|1.0|0.0|RT @jancarlobg: F*ck Donald Trump 
alpha_joe86|Things4Guys|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
alpha_joe86|twitter|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
heyprofbow|iglvzx|0.5766|0.077|0.734|0.189|RT @iglvzx: LMAO. Trump's official website has a glaring XSS vulnerability. You can write in any text to the header.  https://t.co/Ef6oRBK
heyprofbow|t|0.5766|0.077|0.734|0.189|RT @iglvzx: LMAO. Trump's official website has a glaring XSS vulnerability. You can write in any text to the header.  https://t.co/Ef6oRBK
cesarleeon1|Pasion_Basket|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
cesarleeon1|twitter|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
sergiocancelo|Pasion_Basket|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
sergiocancelo|twitter|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
johnathon420|YouTube|0.4404|0.0|0.838|0.162|Ultimate Donald Trump Thug Life Compilation | Funny videos 2016 https://t.co/xi5t4B6tb9 via @YouTube seconds ago  #Trump2016 #TrumpTrain
johnathon420|youtube|0.4404|0.0|0.838|0.162|Ultimate Donald Trump Thug Life Compilation | Funny videos 2016 https://t.co/xi5t4B6tb9 via @YouTube seconds ago  #Trump2016 #TrumpTrain
everydaydolans|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
babybookay|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
babybookay|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Rayaa001|PoppinAssMia|-0.4023|0.311|0.689|0.0|RT @PoppinAssMia: I don't trust Hillary or Trump 
erickd8a|AlecMacGillis|0.0|0.0|1.0|0.0|"RT @AlecMacGillis: All the Trump voters I spoke w/ in PA dismissed his billion-$$ tax writeoff as ""they all do it."" Such a stark example of"
JacobByk|journalsentinel|0.0|0.0|1.0|0.0|"RT @journalsentinel: Preliminary exit polling shows a ""vast gulf of attitudes"" between Trump and Clinton voters in Wisconsin https://t.co/8"
JacobByk|twitter|0.0|0.0|1.0|0.0|"RT @journalsentinel: Preliminary exit polling shows a ""vast gulf of attitudes"" between Trump and Clinton voters in Wisconsin https://t.co/8"
_solleb|FreddieCampion|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
_solleb|twitter|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
lonjoana14|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
lonjoana14|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
heeidi___|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
heeidi___|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
_bombshell_syd|kayla_bayla13|-0.3182|0.315|0.685|0.0|RT @kayla_bayla13: Donald Trump lost https://t.co/7IrlqwgBZ5
_bombshell_syd|twitter|-0.3182|0.315|0.685|0.0|RT @kayla_bayla13: Donald Trump lost https://t.co/7IrlqwgBZ5
gerry_dankowski|PrisonPlanet|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
gerry_dankowski|pittsburgh|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
buffaloon|po_st|-0.2732|0.189|0.811|0.0|Donald Trump Is Suing All The Mexicans https://t.co/GM4XP13b1W via @po_st
buffaloon|wonkette|-0.2732|0.189|0.811|0.0|Donald Trump Is Suing All The Mexicans https://t.co/GM4XP13b1W via @po_st
keepsimpin|Sofy1202|0.5719|0.0|0.748|0.252|RT @Sofy1202: if Trump wins I'll PayPal everyone $1 that RTs this.
madinnz|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
m_skeez|PzFee|-0.7213|0.201|0.799|0.0|RT @PzFee: BREAKING NEWS: TRUMP ASSASSINATED AT RALLY IN OHIO HE HAS BEEN CONFIRMED DEAD. FOLLOW US FOR MORE UPDATES https://t.co/gRNolji43g
m_skeez|twitter|-0.7213|0.201|0.799|0.0|RT @PzFee: BREAKING NEWS: TRUMP ASSASSINATED AT RALLY IN OHIO HE HAS BEEN CONFIRMED DEAD. FOLLOW US FOR MORE UPDATES https://t.co/gRNolji43g
_s0ire|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_s0ire|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
psliker|LOLGOP|0.0516|0.138|0.714|0.148|RT @LOLGOP: EXIT POLL: 3 in 10 Trump supporters had trouble finding the exit to the polls.
BrendanMarks|twitter|0.4767|0.115|0.622|0.263|"Same model says if Trump wins Florida, his chances shoot up to 59%. #ElectionNight #SwingState https://t.co/gDHeVEyxeS"
ang1348|realDonaldTrump|0.0|0.0|1.0|0.0|@realDonaldTrump trump 2016!!
WoodworthElect|SarahPalinUSA|0.0|0.0|1.0|0.0|@SarahPalinUSA My son and I voted for Trump so we can preserve our 2nd Amendment! https://t.co/5QVi2dbKLn
WoodworthElect|twitter|0.0|0.0|1.0|0.0|@SarahPalinUSA My son and I voted for Trump so we can preserve our 2nd Amendment! https://t.co/5QVi2dbKLn
mennahamed8|TheAdly|-0.1027|0.065|0.935|0.0|"RT @TheAdly: #Hillary or #Trump, America will make history today. Either the first female president, or the first mentally challenged one."
SeanKD|SandraTXAS|0.4019|0.057|0.806|0.137|RT @SandraTXAS: Just another good reason #voted #Trump #ElectionDay Bye Bye Amy Schumer will leave if Trump elected https://t.co/SR3Egm
SeanKD|t|0.4019|0.057|0.806|0.137|RT @SandraTXAS: Just another good reason #voted #Trump #ElectionDay Bye Bye Amy Schumer will leave if Trump elected https://t.co/SR3Egm
LMSNCUS|DrMartyFox|-0.0173|0.131|0.741|0.128|RT @DrMartyFox: This Election Is NOT A Choice Between The Lesser Of Two Evils This Is A Choice Between GOOD &amp; PURE EVIL#Voted #Trump On
SinisterCC|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
BDBOY55|DCExaminer|-0.2023|0.121|0.805|0.075|"Voto secreto Trump? Most Hispanics back deportation, want immigration cap cut in half https://t.co/Nje0xALsGV via @DCExaminer"
BDBOY55|washingtonexaminer|-0.2023|0.121|0.805|0.075|"Voto secreto Trump? Most Hispanics back deportation, want immigration cap cut in half https://t.co/Nje0xALsGV via @DCExaminer"
ShrekLover6969|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
LaBar1992|KeithOlbermann|0.0|0.0|1.0|0.0|"RT @KeithOlbermann: Phony ""assassination"" story; FBI; undocumented Melania. The stretch run proved - it's all another Effing Trump Lie http"
BradTurner39|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
jimmymackc|lauraolson|0.0|0.0|1.0|0.0|RT @lauraolson: Pat Toomey says he voted for Donald Trump. #lvelection
BelindaSpeight2|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump now leading IN by 45 points.  RCP has him by 10.  Something is happening.
littleone_96|DaniellBautista|-0.6408|0.458|0.542|0.0|RT @DaniellBautista: FUCK DONALD TRUMP https://t.co/0TUaRyRjgJ
littleone_96|twitter|-0.6408|0.458|0.542|0.0|RT @DaniellBautista: FUCK DONALD TRUMP https://t.co/0TUaRyRjgJ
mmbmak1463|TrumpRising22|0.0|0.0|1.0|0.0|"RT @TrumpRising22: TRUMP - 149,808CLINTON - 62,250"
Miss_TiaJenea|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
williamstubbs95|FunnyPicsDepot|0.3612|0.082|0.781|0.138|RT @FunnyPicsDepot: Stop saying if trump wins yall moving out of the country. Stfu yall cant even move outta ya mommas house https://t
williamstubbs95||0.3612|0.082|0.781|0.138|RT @FunnyPicsDepot: Stop saying if trump wins yall moving out of the country. Stfu yall cant even move outta ya mommas house https://t
alvarezmiguel03|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
alvarezmiguel03|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
_lizcallejas|flawedfacade|0.0|0.0|1.0|0.0|RT @flawedfacade: Y'all talmbout a Trump presidency turning the clock back 500 years when in reality it'll turn the clock back less than 50
Ayoobray_|GIRLHEFUNNY|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
Ayoobray_|twitter|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
femukraine|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
femukraine|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Adriana_Lopez87|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
Adriana_Lopez87|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
hopesprings46|speechboy71|-0.5106|0.202|0.798|0.0|RT @speechboy71: If only Trump had insulted the spouses of every Republican #whatcouldhavebeen https://t.co/ElY8QxJL3U
hopesprings46|twitter|-0.5106|0.202|0.798|0.0|RT @speechboy71: If only Trump had insulted the spouses of every Republican #whatcouldhavebeen https://t.co/ElY8QxJL3U
vviiccttoorr10|ditzkoff|0.0|0.0|1.0|0.0|RT @ditzkoff: Eric Trump gonna Eric Trump https://t.co/JaM3KMhLkL
vviiccttoorr10|twitter|0.0|0.0|1.0|0.0|RT @ditzkoff: Eric Trump gonna Eric Trump https://t.co/JaM3KMhLkL
Adeline_Garrett|YURlPlRATE|0.6633|0.0|0.783|0.217|RT @YURlPlRATE: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
stirlospace|_alastair|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
stirlospace|t|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
gaabiwalsh|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
OnufrijKiselyov|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
OnufrijKiselyov|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
zaylonkitts|EmilyBett|0.0|0.0|1.0|0.0|@EmilyBett TRUMP!!!
xKohai|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
xKohai|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
PantsuitEnFuego|farrightgregy|0.0|0.0|1.0|0.0|"RT @farrightgregy: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
Kofi_ohZmaHn|YemisiSL|0.8555|0.0|0.615|0.385|RT @YemisiSL: I actually don't understand black people that support Trump. Like I'd love to ask a few questions. Forreal
ctconnolly56|TeresaEdelglass|0.4019|0.0|0.838|0.162|RT @TeresaEdelglass: #Trump's African-American Support Highest For #GOP Since 1960 #VoteTrump #BlackVote #Trump2016 #AmericaFirst #MAGA h
MericanDude|Breaking911|0.0|0.0|1.0|0.0|RT @Breaking911: Trump Voters Claiming Ballots Defaulting To Clinton https://t.co/tNSlrPtv8F
MericanDude|breaking911|0.0|0.0|1.0|0.0|RT @Breaking911: Trump Voters Claiming Ballots Defaulting To Clinton https://t.co/tNSlrPtv8F
JazmineMejia14|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
JazmineMejia14|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
ReviewDuckUSA|bigmates|0.0|0.0|1.0|0.0|@bigmates trump
3arbylka|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
3arbylka|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
kirstenstauffe1|LondraPolitics|0.0|0.0|1.0|0.0|"RT @LondraPolitics: According to the Turkish media funded by Erdogan, here is the first #ElectionNight exit poll results;Hillary: 20%Tru"
jsrroger|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @Slate @votecastr @LilSteelerGirl @DebAlwaystrump @Kerri1111 TRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLID
britnaaymariie|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
britnaaymariie|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
MarkGreen88|matt_dederer|-0.4023|0.153|0.847|0.0|RT @matt_dederer: When you don't trust your own wife to vote for you #Trump #electionday https://t.co/7oNK4EmijQ
MarkGreen88|twitter|-0.4023|0.153|0.847|0.0|RT @matt_dederer: When you don't trust your own wife to vote for you #Trump #electionday https://t.co/7oNK4EmijQ
ftvoc|R5Eileen|0.8398|0.104|0.347|0.549|"RT @R5Eileen: Please God, let Trump be the clear cut winner! https://t.co/XE5Gs3UXEA"
ftvoc|twitter|0.8398|0.104|0.347|0.549|"RT @R5Eileen: Please God, let Trump be the clear cut winner! https://t.co/XE5Gs3UXEA"
CCrusherP|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
sirdrano|PerlinaCucina|0.296|0.0|0.891|0.109|RT @PerlinaCucina: I voted for Donald Trump and Mike Pence. Will you join me? Find your polling place: https://t.co/W0iumzOnqn #TrumpTrain
sirdrano|vote|0.296|0.0|0.891|0.109|RT @PerlinaCucina: I voted for Donald Trump and Mike Pence. Will you join me? Find your polling place: https://t.co/W0iumzOnqn #TrumpTrain
supbrea|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Blonde_Politico|fmlannalisa|0.3612|0.0|0.878|0.122|@fmlannalisa because I'm not voting with my vagina.  Sounds like you need a gynecologist and not a president.  #MAGA #Election2016 #Trump
heatcost245780|megynkelly|0.0|0.0|1.0|0.0|"RT @megynkelly: 18 electoral votes are up for grabs in #Ohio, and the states own Republican Gov. John Kasich says he did not vote for #Tru"
JakaylaLovesYou|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
JakaylaLovesYou|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
TrumpWithUSA|Democrat_4Trump|0.5106|0.062|0.782|0.156|"RT @Democrat_4Trump: CNN CAUGHT: Blitzer talks, CNN flashes a Trump Florida win for 2 seconds then takes it offline quick. Why don't they s"
andysRoses|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
KaylaSpriggs|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
AngelNapoles4|_Makada_|0.0|0.0|1.0|0.0|RT @_Makada_: I #voted for Donald Trump for POTUS! AMERICA FIRST! #ElectionDay https://t.co/eQuXYsXvg9
AngelNapoles4|twitter|0.0|0.0|1.0|0.0|RT @_Makada_: I #voted for Donald Trump for POTUS! AMERICA FIRST! #ElectionDay https://t.co/eQuXYsXvg9
kLodeserto|theglobaluniter|0.0|0.0|1.0|0.0|RT @theglobaluniter: If you live in the Panhandle area of Florida we need you to go and #Vote #Trump.A call to action by .@DonaldJTrumpJ
tanner_coleman|jasonvolack|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
tanner_coleman|twitter|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
murphyj21|surfermom77|0.0|0.0|1.0|0.0|"RT @surfermom77: Twitter &amp; FB R begin inundated wt reports of Elec.fraud, voting irregularities &amp; discrimination against Trump Votershttps"
fruace|oneofonealbum|0.5719|0.0|0.821|0.179|RT @oneofonealbum: If Trump   Wins The Election I Am Moving   Out Of The Country  Goodbye   America   Hello   SHINee Wo
WagnerJwagner23|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
VonWally|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
EEGRC98|0hour|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
EEGRC98|twitter|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
charley_ck14|hipsterocracy|0.5719|0.0|0.764|0.236|"RT @hipsterocracy: If Trump somehow wins, Golden Corral is gonna be lit tonight."
gutierrezy14|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
gutierrezy14|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
HmartinPalm|Koxinga8|0.6174|0.053|0.758|0.189|RT @Koxinga8: Start Packing &amp; Booking Removalist Yet???  16 Celebrities Who Will Leave the U.S. if Trump Wins  https://t.co/RXTDdiav1Q
HmartinPalm|breitbart|0.6174|0.053|0.758|0.189|RT @Koxinga8: Start Packing &amp; Booking Removalist Yet???  16 Celebrities Who Will Leave the U.S. if Trump Wins  https://t.co/RXTDdiav1Q
ceciliagomezsa|Gloful_|-0.6486|0.301|0.699|0.0|RT @Gloful_: If you voted for Donald trump ya moms a whore
silverfoxmedia1|mitchellvii|0.34|0.0|0.893|0.107|"RT @mitchellvii: I expect Trump to win KY and IN, but not by 50 points.  We'll see if anything near that holds."
goodyk|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
FACT_gr|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
FACT_gr|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
VonFuzzyhead|cliffschecter|0.2263|0.0|0.921|0.079|"RT @cliffschecter: In Clarke Cnty Nevada, Trump sues 2 throw out votes. In Durham, Ds sue to allow more ppl 2 vote. Any questions? https://"
VonFuzzyhead||0.2263|0.0|0.921|0.079|"RT @cliffschecter: In Clarke Cnty Nevada, Trump sues 2 throw out votes. In Durham, Ds sue to allow more ppl 2 vote. Any questions? https://"
felipe_lab|twitter|0.5719|0.137|0.497|0.366|So far Kentucky n Indiana Trump supposed to win. No surprise https://t.co/I6u4WdzPZH
Redjen40J|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
JankowiakJoAnn|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
JankowiakJoAnn|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
svogel2|movement_trump|0.6689|0.0|0.793|0.207|"RT @movement_trump: Do you really want another flaming liberal on the Supreme Court?  If not, you must vote for Donald J Trump TODAY! https"
CopeGerry|LeafyIsHere|0.4238|0.139|0.589|0.272|"RT @LeafyIsHere: If Trump wins I'll release nudes, not a joke"
MCRWillCarryOn_|BoofBaldy|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
MCRWillCarryOn_|twitter|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
derya555|AdamsFlaFan|0.0|0.0|1.0|0.0|"RT @AdamsFlaFan: Donald Trump 'needs a test of his sanity,' says 105-year-old voter https://t.co/4nLgHbGy2x"
derya555|newsweek|0.0|0.0|1.0|0.0|"RT @AdamsFlaFan: Donald Trump 'needs a test of his sanity,' says 105-year-old voter https://t.co/4nLgHbGy2x"
kiraaaax3_|BeenBabyKi|0.3612|0.0|0.8|0.2|RT @BeenBabyKi: Not Voting At All Is Like Voting For Trump
cguerra121|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
BMGConsulting|instagram|0.5411|0.0|0.589|0.411|Vote Trump to save America! https://t.co/4WW0EeZEvO
deltarag14|damaninthearena|0.0|0.0|1.0|0.0|RT @damaninthearena: @Vendetta92429 @antimarxis_ this map is BS!! I'm in southern Cali and in a line of 50+ people; Black White Hispanic As
sheryl_harvey|Cory_1077|0.0|0.0|1.0|0.0|RT @Cory_1077: VOTE TRUMP To get rid if the #PoliticalCorruption in our Country #MakeAmericaGreatAgain   #MakeAmer
be_emb|twitter|0.0|0.0|1.0|0.0|#FoxNews2016 My 18 year old daughters first vote. Go Trump!! https://t.co/v5AoHQc7kg
KeithZ07|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
xkr99|GartrellLinda|0.2714|0.0|0.905|0.095|RT @GartrellLinda: Important! RTGET OUT THERE &amp; VOTE TRUMPSTERSVERY TIGHT in Florida panhandle. Call everyone you know to get those Trump
bobnfn1|TheDonaldNews|-0.783|0.346|0.654|0.0|@TheDonaldNews @ed_hooley @realDonaldTrump @DanScavino @Always_Trump Keep voting!! We need to crush these evil people! #DrainTheSwamp
USAHipster|WDFx2EU8|0.0|0.0|1.0|0.0|"RT @WDFx2EU8: BOOM: 94 y.o. lady in line, Votes TRUMP, last time she voted...was Franklin Roosevelt! #electionday"
greigo_uk|Miserable_Me1|0.5622|0.0|0.623|0.377|@Miserable_Me1 HOPE ITS NOT TRUMP FACE THO
tothemaxxi|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
tothemaxxi|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
WD_Lady|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
WD_Lady|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
BegiiiGiles|pharris830|-0.5719|0.209|0.791|0.0|RT @pharris830: Furious Trump Fans Just Found Out They Have To Register To Vote - https://t.co/qgV2c1svBf
BegiiiGiles|occupydemocrats|-0.5719|0.209|0.791|0.0|RT @pharris830: Furious Trump Fans Just Found Out They Have To Register To Vote - https://t.co/qgV2c1svBf
kevole|instagram|0.0|0.0|1.0|0.0|The polls are about to close.#getyourpopcornready #electionnight #Trump #clinton https://t.co/hpio9fRlGG
fflooff|NathanZed|0.5719|0.0|0.866|0.134|RT @NathanZed: if trump wins im moving to my grandmas house. she still live in america this don't got anything to do with politics I just m
paigeneely4|b0rby|0.0|0.0|1.0|0.0|RT @b0rby: Thoughts on Trump https://t.co/1KWxB5ciHT
paigeneely4|twitter|0.0|0.0|1.0|0.0|RT @b0rby: Thoughts on Trump https://t.co/1KWxB5ciHT
ASauer65|EntheosShines|0.4404|0.0|0.861|0.139|RT @EntheosShines: @iamgavinjames A Gift To You - The Trump Movement Video Storybook Of Past 18 Months @DanScavino @Harlan @Cernovich https
streetwise_IT|DanScavino|0.0|0.0|1.0|0.0|RT @DanScavino: Trump Campaign Headquarters-'TOP CANDIDATE QUALITY: CAN BRING CHANGE:TRUMP: 82%CLINTON: 13%#iVoted #ElectionNight #MAGA
tdobbs431|twitter|0.6486|0.0|0.569|0.431|"Thank,you Mr.Trump for giving American a voice again n hope https://t.co/ctEfNLhcds"
darby__ann|twitter|-0.34|0.272|0.543|0.185|"A whole lot a ignorance in one little girl. I'm a trump supporter, no one is useless. Honestly honey, you need so e https://t.co/4gLG1O2Q4F"
frespirit01|MagicRoyalty|0.8225|0.0|0.714|0.286|RT @MagicRoyalty: WOW: another proof of #VoterFraud!! Machine refuses to allow vote for Trump!!RT b/c Media will never report this! http
_NoFilter_|_ShowNoLovee|0.0|0.0|1.0|0.0|@_ShowNoLovee trump and Hillary 
VeeLo_Greene|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
Kinjo_Goldbar|mitchellvii|0.4404|0.0|0.805|0.195|"RT @mitchellvii: Trump leads IND 72-25.  Good Lord people, something is happening here."
gibsonnbecca|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
gibsonnbecca|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
kathyfisher10|JMilesColeman|0.0|0.0|1.0|0.0|RT @JMilesColeman: Elliott County KY going 66% for Trump. This is probly the year it finally buckles to the Rs. #kyvote
HookerBot5000|farrell_nic|-0.2023|0.096|0.904|0.0|Sobering midnight (GMT) text from @farrell_nic : 'WHAT IF WE WAKE UP AND TRUMP IS PRESIDENT'. I can't sleep now 
Brendalea414|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
s_hutchy|Felangomango|0.4404|0.0|0.734|0.266|RT @Felangomango: Good Morning to everyone except Donald Trump
IM_extrAVAgant|Inc|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
IM_extrAVAgant|t|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
kathicolorado|marshawright|0.0|0.0|1.0|0.0|RT @marshawright: KENTUCKY EARLY RESULTS EXIT POLLSEARLY LEADS: POTUS ALERTTRUMP 72.7%CLINTON 24.6%#ElectionNight #electionday #IVOTE
saveAmerica123|enfingercolton2|0.3802|0.0|0.776|0.224|@enfingercolton2 Please consider this article before voting for Trump! https://t.co/3D6lxGFB5v
saveAmerica123|medium|0.3802|0.0|0.776|0.224|@enfingercolton2 Please consider this article before voting for Trump! https://t.co/3D6lxGFB5v
LeDeplorables|WDFx2EU8|0.8443|0.0|0.597|0.403|"RT @WDFx2EU8:  BREAKING: WOW!!! At the last minute, Chris Matthews endorses #Trump!!! #ElectionDay  https://t.co/FjeNWIsACt"
LeDeplorables|twitter|0.8443|0.0|0.597|0.403|"RT @WDFx2EU8:  BREAKING: WOW!!! At the last minute, Chris Matthews endorses #Trump!!! #ElectionDay  https://t.co/FjeNWIsACt"
DrunkyBorghy|twitter|0.0|0.0|1.0|0.0|#Election2016 NOT DONALD TRUMP NOT DONALD TRUMP NOT DONALD TRUMP https://t.co/VbiTfZ2yYX
bearoserod|BuzzFeedNews|-0.7028|0.271|0.729|0.0|"RT @BuzzFeedNews: 29 Most WTF Moments Of The Election: Hillary's Trump ""Joke"" #ElectionDay https://t.co/PNF7xkBxgB"
bearoserod|twitter|-0.7028|0.271|0.729|0.0|"RT @BuzzFeedNews: 29 Most WTF Moments Of The Election: Hillary's Trump ""Joke"" #ElectionDay https://t.co/PNF7xkBxgB"
AntonLaGuardia|khalafroula|0.7506|0.0|0.701|0.299|"RT @khalafroula: Looks like Trump got his wall after all. A wall of beautiful voters, Latinos in nevadahttps://t.co/ar83t8XqUx"
LivingBigly|Thomas1774Paine|-0.2023|0.087|0.913|0.0|RT @Thomas1774Paine: Notice you never see #Clinton voters complaining the voting machine changed their vote to #Trump? Wonder why ...
votingtrump|NYtoKYChristian|0.0|0.0|1.0|0.0|"RT @NYtoKYChristian: @bitsy423 @cnoss53 @zclove2bme @dkarnok Long Island NY Hundreds in pro-Trump parade shouting ""lock her up!"" #votedTrum"
toddage_cheese|mlissa1|-0.2263|0.142|0.751|0.107|RT @mlissa1: I am a Mexican American that lives in South Texas. Unlike Ana Navarro I clearly heard when Trump said Illegal immigrants. I vo
Haley_Greentree|Thomas1774Paine|0.0|0.0|1.0|0.0|RT @Thomas1774Paine: Female #Trump voter hammers CNN. Yinz shouldn't have asked the question if Yinz at CNN didn't know the answer. Google
simonstanton|instagram|0.0|0.0|1.0|0.0|"At work, reviewing analytics language breakdown, this appears. Vote trump??? google googleanalytics https://t.co/TGSYsqumHg"
rlgordon18_ruth|FrankLuntz|0.25|0.0|0.889|0.111|RT @FrankLuntz: BREAKING: Watch Michigan.Working-class turnout is looking much higher than expected. Trump may actually have a chance.  #
jim_hollifield|FrankLuntz|-0.1027|0.055|0.945|0.0|RT @FrankLuntz: The turnout in Democratic Philadelphia is so high that it's hard to see Trump overcoming it in the rest of the state.  #Ele
Katiecook55|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
Katiecook55|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
blessedboymama|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: We don't know the following:1) How many Democrats are voting Trump.2) How many Independents are voting Trump.Relax.
Quany_Flamez|ItsChinaa_|0.0|0.0|1.0|0.0|RT @ItsChinaa_: If donald trump gets elected as president.. 9/10 he will get impeached.
DeadlineDavis|anthonyalsop|-0.4215|0.286|0.714|0.0|"@anthonyalsop ""Trump cheats vote and makes it informal"""
DONNABELLINI1|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
DONNABELLINI1|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
Skydawgy1|TomiLahren|0.4717|0.0|0.861|0.139|RT @TomiLahren: If you're not voting for Trump don't you dare bitch when we get Hillary. Real talk. #MAGA #ElectionDay
USA_with_Trump|jackbgoode1|0.6249|0.0|0.728|0.272|RT @jackbgoode1: Great question  - VOTE TRUMP @DonaldTrumpVote @USFreedomArmy @Karennola719 @Jnbarke @realDonaldTrump https://t.co/O3B8mIkz
USA_with_Trump|t|0.6249|0.0|0.728|0.272|RT @jackbgoode1: Great question  - VOTE TRUMP @DonaldTrumpVote @USFreedomArmy @Karennola719 @Jnbarke @realDonaldTrump https://t.co/O3B8mIkz
lmvanness|majtague|0.0|0.0|1.0|0.0|"RT @majtague: #DistractMeWithAnElectionPoemRoses are red,Trump's out there hatin' But if you vote we can say: https://t.co/0Mi3dsthp9"
lmvanness|twitter|0.0|0.0|1.0|0.0|"RT @majtague: #DistractMeWithAnElectionPoemRoses are red,Trump's out there hatin' But if you vote we can say: https://t.co/0Mi3dsthp9"
MaximAlesandr|Reevellp|0.4019|0.0|0.881|0.119|RT @Reevellp: In #Moscow there is a Trump party in-full swing- pro-Kremlin activists gathered in a bar for the results. Giant portrait of T
ToeKnee2GX|AceHudsonJr|0.4404|0.0|0.775|0.225|@AceHudsonJr @jhood102 SMFH hope Trump gets elected so u can be deported
WryghtSparrow|BREAKING_PTV|0.0|0.0|1.0|0.0|"RT @BREAKING_PTV: Early results: Trump leads Clinton in states of Indiana, Kentucky, new Hampshire#ElectionDay #Election2016 https://t.co"
WryghtSparrow|t|0.0|0.0|1.0|0.0|"RT @BREAKING_PTV: Early results: Trump leads Clinton in states of Indiana, Kentucky, new Hampshire#ElectionDay #Election2016 https://t.co"
jtmcewan11|Nija315|0.2185|0.192|0.533|0.275|RT @Nija315: Donald trump is winning the popular vote... SHIT IS ABOUT TO GET REAL
HazelOsterhout|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Running_creek|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
siaayrom|ananavarro|-0.2732|0.087|0.913|0.0|"RT @ananavarro: Hey Nevadans, u know why Trump is suing? To keep Hispanics from polls b/c he knows we're voting against him. Redouble your"
Nise_Renee|dwontlose|-0.25|0.366|0.323|0.312|RT @dwontlose: Trump supporters are truly dumb as fuck https://t.co/xblDZE2RcA
Nise_Renee|twitter|-0.25|0.366|0.323|0.312|RT @dwontlose: Trump supporters are truly dumb as fuck https://t.co/xblDZE2RcA
pau2la057328721|manusartorius02|-0.6408|0.514|0.486|0.0|RT @manusartorius02: FUCK OFF TRUMP 
russmove|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
zapoteco|xeni|-0.6369|0.257|0.743|0.0|"RT @xeni: From our archives: Donald Trump confirms, then denies, his father's arrest at a KKK rally https://t.co/JvIzuUcE5h"
zapoteco|boingboing|-0.6369|0.257|0.743|0.0|"RT @xeni: From our archives: Donald Trump confirms, then denies, his father's arrest at a KKK rally https://t.co/JvIzuUcE5h"
TheNoahBrinson|Patterrz|-0.1336|0.296|0.704|0.0|RT @Patterrz: Serious tho don't elect Trump pls
jesssica_z|twitter|0.6486|0.091|0.588|0.321|This has got to be a joke you CAN NOT seriously let trump win https://t.co/HIx0dsmMva
DlCKFORD|Miikeyyv|0.0|0.0|1.0|0.0|@Miikeyyv @ggullotti1 @jojo_bear32 @jackwilsonnnnnn still don't see connection to trump
bringitbri_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
GagAlexFrance|musicnews_facts|0.4404|0.0|0.873|0.127|"RT @musicnews_facts: Trump supporters are calling out Hillary Clinton and Lady Gaga for wearing this ""Nazi Hitler"" uniform... When it's Mic"
BrianMyrieSalsa|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
BrianMyrieSalsa|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
newsbreak|cnn|0.0|0.0|1.0|0.0|#cnn First returns: Trump leads in Indiana https://t.co/oerqDOZJnL
SOgnenis|roweafr|0.5859|0.0|0.612|0.388|RT @roweafr: the joy #TRUMP #USElection2016 https://t.co/2RwskxNZYk
SOgnenis|twitter|0.5859|0.0|0.612|0.388|RT @roweafr: the joy #TRUMP #USElection2016 https://t.co/2RwskxNZYk
aamilgerard|NathanZed|0.5719|0.0|0.866|0.134|RT @NathanZed: if trump wins im moving to my grandmas house. she still live in america this don't got anything to do with politics I just m
TheEfbe|WhoadieBrees|-0.4003|0.152|0.848|0.0|RT @WhoadieBrees: Niggas with white gfs RT @lovemeGabbi: Who is this 8% voting for trump?! https://t.co/qsNsQ3stvV
TheEfbe|twitter|-0.4003|0.152|0.848|0.0|RT @WhoadieBrees: Niggas with white gfs RT @lovemeGabbi: Who is this 8% voting for trump?! https://t.co/qsNsQ3stvV
JVjett|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
estefanigarciaO|richchigga|0.3182|0.0|0.85|0.15|RT @richchigga: please do not vote for donald trump so i can come to america
jdashstylez|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
jdashstylez|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
realevie_|lovelykmx|-0.3724|0.358|0.466|0.177|RT @lovelykmx: Trump can't seriously win
itvnews|twitter|-0.7351|0.307|0.693|0.0|Jesse Jackson says US has ideological struggle similar to that of America's civil war #Election2016 https://t.co/QMIpmJTe40
BillLonbeck|mitchellvii|0.3182|0.0|0.723|0.277|RT @mitchellvii: Trump leads Kentucky 77-20. :-)
MrGlennoo|MerlotGrey|-0.296|0.115|0.885|0.0|RT @MerlotGrey: @reeeaaalllyreal @mitchellvii Stop posting bs.  CNN is not privy to the internals of the Trump camp.
vhfancc|CatalenaNikole|-0.4215|0.241|0.62|0.139|"@CatalenaNikole @8simon9 Now thats a real USA lover , man on the verge of death still fights to cast ballot for Trump ."
my_eskie|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
my_eskie|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
jbritta|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
KonorFelix|troyesivan|-0.3182|0.133|0.867|0.0|RT @troyesivan: i dont mean to be a tease but....like...imagine not having to hear about donald trump anymore 
buckitman|michaelharrisdr|0.4404|0.0|0.805|0.195|"RT @michaelharrisdr: #TrumpWinsBecause  says Patriots' Tom #Brady, Bill #Belichick supporting him @CNNPolitics https://t.co/kCFsGmSkPc"
buckitman|edition|0.4404|0.0|0.805|0.195|"RT @michaelharrisdr: #TrumpWinsBecause  says Patriots' Tom #Brady, Bill #Belichick supporting him @CNNPolitics https://t.co/kCFsGmSkPc"
susan_250|BiccyM|-0.7579|0.246|0.754|0.0|RT @BiccyM: I know it is lazy to assume all Trump fans are stupid but there is a deep rooted educational problem that has allowed him to ge
naeebrazy|iam_dezziedoll|0.0|0.0|1.0|0.0|RT @iam_dezziedoll: If you voted for Donald trump and you black bye you white now 
bigchetti|40oz_VAN|0.5719|0.0|0.821|0.179|RT @40oz_VAN: How are you leaving the country if Trump wins if you've never even left your city?
SandraKennett1|LouDobbs|-0.7574|0.372|0.544|0.083|"@LouDobbs Hillary isn't well liked by people, while Donald Trump is loved by people, but not well liked by the biased MSM."
MeganNemec|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
MeganNemec|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
RickyFoley|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
RickyFoley|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
thisboijesse|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
tynmadimom|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: RCP average in Indiana has Trump up 10.  He is currently up close to 50!!!  Monster vote?  Crossovers?
SomeGuysCat|JohnFromCranber|0.6739|0.0|0.835|0.165|RT @JohnFromCranber: It's All About Turnout. Typically Only About 1/2 Vote. If All the Folks who Prefer Trump Over Hillary Vote - WE WIN IN
Humdingerding|NRO|0.0|0.0|1.0|0.0|"RT @NRO: Early Exit Polls: Trump Opens YUGE Gap between College-Educated, Non-College-Educated Whiteshttps://t.co/ADpCNhYfiC #ElectionNight"
Trump_45th_Pres|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: Your vote right now is more than just the next 4 years. It is a generational vote. One that will be felt for decades. #
vekmar|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
chinosanap|timinhoustontex|0.0|0.0|1.0|0.0|RT @timinhoustontex: #TrumpTrain #NAACP #msnbc #cnn #ImWithHer #NYTimes #foxnews #bikers4trump #cnbc #abc #loudobbs All of us must ge
spiritofshiloh|staffsgtshawnb2|0.5267|0.0|0.726|0.274|RT @staffsgtshawnb2: #FoxNews2016.  trump is winning new Hampshire. 52 41
SandyKuti|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: Right now, Trump is making up more than half of Obama's entire 2012 margin of victory in FL in JUST ONE COUNTY!"
MrBrownThumb|twitter|-0.4588|0.13|0.87|0.0|"If you're not voting 'cause the lines are too long, just imagine the lines for forced labor and deportation camps u https://t.co/5ekqXTvE3i"
TheAmishDude|AG_Conservative|-0.3612|0.172|0.712|0.116|"RT @AG_Conservative: Again, Trump now only guaranteed ""amnesty,"" but also made border security unpopular. He hurt every cause he claimed to"
whateverlyss|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
whateverlyss|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
kvnax|l4444k|0.0|0.0|1.0|0.0|RT @l4444k: Snoop Dogg @ Donald Trump Roast https://t.co/SkVuien0t8
kvnax|twitter|0.0|0.0|1.0|0.0|RT @l4444k: Snoop Dogg @ Donald Trump Roast https://t.co/SkVuien0t8
sassyfairex|caramelthot|-0.1655|0.064|0.936|0.0|"RT @caramelthot: my neighbor just told me someone stole her trump sign last night &amp; i acted all shocked, but little does she know i was the"
miatorch|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
miatorch|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
DotCalm_6|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
haddynuff|StopStopHillary|0.0|0.0|1.0|0.0|RT @StopStopHillary: FIRST POLLS FOR KENTUCKY TRUMP 78%HILLARY 18%
ARepublic|KellyannePolls|0.7096|0.0|0.781|0.219|RT @KellyannePolls: Trump Campaign &amp; RNC @Reince hand in glove. This is about GOP elected officials bragging they voted 3rd party or skippe
7Canyons|Cernovich|0.0|0.0|1.0|0.0|RT @Cernovich: Two votes for Trump on #ElectionDay!#MAGASelfie https://t.co/nOtQqiSW36
7Canyons|twitter|0.0|0.0|1.0|0.0|RT @Cernovich: Two votes for Trump on #ElectionDay!#MAGASelfie https://t.co/nOtQqiSW36
sumbodysbabygrl|letters2donald|-0.5255|0.145|0.855|0.0|"RT @letters2donald: Children's letters to Donald Trump:  Some of your fans lie even worse than you do. I bet that's a relief!Connor F., a"
kristinkgl|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
kristinkgl|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
ChandracCl|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Ptmurf1016|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
iChristNews|christianitytoday|0.2023|0.0|0.878|0.122|Top 10 Stats Explaining the Evangelical Vote for Trump or Clinton https://t.co/4jQc5fZEdq #Christian #News
aislam_|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
cairnstoon|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
cairnstoon|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
laurenalexis26|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
laurenalexis26|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
Donatopanic|DonaldJTrumpJr|0.8442|0.0|0.435|0.565|@DonaldJTrumpJr @EricTrump god let mr trump win save our country
GreeneRbt|JonahNRO|-0.3612|0.102|0.898|0.0|RT @JonahNRO: 1. Trump is more liberal than Bush. 2. I criticized Bush's liberalism. 3. There are *many* reasons to object to Trump other t
JoeRiggs10|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
lampieeee9|FoxNews|0.6124|0.0|0.778|0.222|@FoxNews we early voted for Trump in Maryland our lovable pit raven sums it up
prof_gabriele|trump_cake|0.0|0.0|1.0|0.0|Guys follow @trump_cake now
srslyfrank|niicest|0.0|0.0|1.0|0.0|"RT @niicest: If you're Hispanic/Latino voting trump, ima need u to write a 10 page essay explaining yo self, so I can then spit on it throw"
caaroliinam|VanityFair|0.4019|0.084|0.756|0.16|RT @VanityFair: Nevada judge becomes hero for telling Trump lawyer to sit down over absurd voter lawsuit https://t.co/Q6ogpd1NNA https://
caaroliinam|vanityfair|0.4019|0.084|0.756|0.16|RT @VanityFair: Nevada judge becomes hero for telling Trump lawyer to sit down over absurd voter lawsuit https://t.co/Q6ogpd1NNA https://
KarlaPa23670577|gothamist|-0.6597|0.375|0.625|0.0|Rebels Beamed Anti-Trump 'Star Wars' Scroll By Darth Trump's Tower https://t.co/pEFyDlJGU0
yomemy|HorridPineapple|0.4404|0.0|0.818|0.182|RT @HorridPineapple: It's how you weed out the trump supporters from your life https://t.co/8fZqzhaJFX
yomemy|twitter|0.4404|0.0|0.818|0.182|RT @HorridPineapple: It's how you weed out the trump supporters from your life https://t.co/8fZqzhaJFX
CPCB|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
CPCB|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
mamasaurusof2|thehill|0.5106|0.0|0.784|0.216|RT @thehill: Early exit poll: Clinton tops Trump in ground game https://t.co/l0AGQ5nhc0 https://t.co/3n0aSSL3kn
mamasaurusof2|thehill|0.5106|0.0|0.784|0.216|RT @thehill: Early exit poll: Clinton tops Trump in ground game https://t.co/l0AGQ5nhc0 https://t.co/3n0aSSL3kn
Sherri1030|mitchellvii|0.5267|0.0|0.673|0.327|RT @mitchellvii: I see Trump winning MI and CO.
AbhayJhaveri|immoumita|0.2263|0.0|0.881|0.119|"RT @immoumita: News channels had prepared for Clinton n trump, Modi came out of syllabus  #currencyswitch"
fergesor|hrtablaze|0.9207|0.0|0.645|0.355|RT @hrtablaze: My Bernie Sanders loving nephew who has been messing with me all election just told me he voted TRUMP !!! WOOT WOOT ! #elect
sameoldsxlena|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
sameoldsxlena|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
Jake_Learned|Bernie_Facts|0.6812|0.0|0.765|0.235|@Bernie_Facts so Trump should win? You realize that's what you're saying? Are you guys even pro-Bernie?
mariaisimoza|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
mariaisimoza|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
andrialisa24|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: I wonder if anyone at Trump campaign is busily looking to see if Nevada Judge has Hispanic ancestry somewhere in her ba
RidesPet|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you voted for TRUMP! #ElectionDay #Vote #Vote2016
bleudawn7|alicebonasio|-0.5423|0.2|0.8|0.0|RT @alicebonasio: Millennials: get off your ass and #VOTEHILLARY NOW https://t.co/VlfdwzM0LX  #ElectionFinalThoughts #Election2016 @qz #br
bleudawn7|qz|-0.5423|0.2|0.8|0.0|RT @alicebonasio: Millennials: get off your ass and #VOTEHILLARY NOW https://t.co/VlfdwzM0LX  #ElectionFinalThoughts #Election2016 @qz #br
spdygdallas|RalstonReports|0.0|0.0|1.0|0.0|"RT @RalstonReports: Trump: ""We have reason to believe too many Dems voted.""Judge: ""But it's the law to let people in line vote.""Trump: ""B"
copstaff|conspiracyoutpost|0.0|0.0|1.0|0.0|NOOOO Waaaaaaaayy!!!!: Clinton | Kaine V Trump | Pence Cain&gt;fenced garden  V  Trumpets https://t.co/DRMWmeSbGX https://t.co/3XvKZjn4Jd
JarrodSHagenman|Variety|-0.8176|0.362|0.638|0.0|@Variety assholes.  That's automatic vote for Trump. Leave it to three #bushes to fuck up an election #imwithher
pewdrdad|youngcons|0.4404|0.0|0.847|0.153|"First Early Exit Polls Just Released, and They Point Towards Good News for Trump https://t.co/9CPoJdWqrG via https://t.co/2ox3KTKlKx"
DawnSwe12515208|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: Folks, if you are at work and trying to decide whether to still vote for Trump,GO VOTE, MAKE HISTORY!"
AshandCinders|kcinderfell|0.5719|0.073|0.664|0.262|RT @kcinderfell: regardless of what happens if you live in the us please be careful because no matter what trump supporters are going to be
DANNYHOAGLAND1|twitter|-0.368|0.336|0.664|0.0|TRUMP TRAIN IS UNSTOPPABLE   - PATTON https://t.co/crSYvgLxQ5
AmberGirl3|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
LavelleGerald|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
LavelleGerald|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
ApocalypticaNow|jesseberney|-0.5267|0.208|0.69|0.102|RT @jesseberney: Trump has broken a lot of norms but I like the new tradition he established that the loser has to eat a cake of himself lo
karaaaMarieee7|brooke7899|0.0|0.0|1.0|0.0|TRUMP 2016 BUILD THAT WALL @brooke7899 https://t.co/ytteudfrwx
karaaaMarieee7|twitter|0.0|0.0|1.0|0.0|TRUMP 2016 BUILD THAT WALL @brooke7899 https://t.co/ytteudfrwx
_Byethai|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_Byethai|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
tkamins123|dmckinney218|0.0|0.0|1.0|0.0|RT @dmckinney218: Hispanics voting for Donald Trump! https://t.co/Uq66TaDVQ2
tkamins123|twitter|0.0|0.0|1.0|0.0|RT @dmckinney218: Hispanics voting for Donald Trump! https://t.co/Uq66TaDVQ2
julieorth2|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
corgilessEmily|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
corgilessEmily|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
miflorhermosa|caramelthot|-0.1655|0.064|0.936|0.0|"RT @caramelthot: my neighbor just told me someone stole her trump sign last night &amp; i acted all shocked, but little does she know i was the"
beltranaminta|lowelljohnsonjr|0.2023|0.0|0.904|0.096|"RT @lowelljohnsonjr: Top story: Some Trump Voters Reporting Ballots Switching To Clinton  CBS Pitts https://t.co/2rVmyqslFQ, see more htt"
beltranaminta|pittsburgh|0.2023|0.0|0.904|0.096|"RT @lowelljohnsonjr: Top story: Some Trump Voters Reporting Ballots Switching To Clinton  CBS Pitts https://t.co/2rVmyqslFQ, see more htt"
bistrogal2|twitter|0.5599|0.0|0.859|0.141|"PLEASE EVERYONE.GET OUT &amp; VOTE FOR TRUMP! EVEN IF YOU HAVE A COLD, APPT - ANY REASON, JUST GET OUT &amp; VOTE! DRAIN TH https://t.co/Z7UKiWzkHL"
tronnorxdosogas|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
Pro_America1776|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
Its_Freddie|lou_snatch|0.5859|0.0|0.612|0.388|RT @lou_snatch: @Its_Freddie trump gonna win bruhh
sharsheepdog|MattGertz|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
sharsheepdog|twitter|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
shxmvllnv|vibeeeez|-0.5574|0.261|0.739|0.0|RT @vibeeeez: prediction: Hillary Clinton is our next present &amp; everyone is shocked Trump lost
FirstNameMiaa|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
FirstNameMiaa|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
jktrails13|BretBaier|-0.1531|0.117|0.789|0.094|GOP not voting Trump is like not getting in the last lifeboat on the Titanic because it's the wrong color. #Election2016 @BretBaier @FoxNews
GoldenPhiliRoll|Aimee_P_R|0.0|0.0|1.0|0.0|RT @Aimee_P_R: Trump isn't allowed to control his own Twitter account but some people think he should control one of the world's most power
mariaeke|bipartisanreport|0.2103|0.0|0.857|0.143|BREAKING: FBI STUNS America With Election Day Trump/Russia Warrant Announcement (DETAILS) https://t.co/MSmf7cvINR
timfromhouston|twitter|0.3612|0.0|0.8|0.2|Arriving on the TL to watch the #trump #meltdown like: https://t.co/VLQOgyCQAh
FrannieC_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
RockieBilbrey|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
RockieBilbrey|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
Deserie_Larios|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
Deserie_Larios|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
shar_veshh|BazK10|0.5719|0.0|0.73|0.27|RT @BazK10: I will eat this if trump wins the election  https://t.co/SGLHSg7MmO
shar_veshh|twitter|0.5719|0.0|0.73|0.27|RT @BazK10: I will eat this if trump wins the election  https://t.co/SGLHSg7MmO
kabbath|KHQA|0.0|0.0|1.0|0.0|RT @KHQA: Eric Trump illegally posts pic of completed NY ballot on Twitterhttps://t.co/o3ic19ZzeU
focused_4|Chico_Mills|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
focused_4|twitter|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
USAgladiator2|smoothkobra|-0.7964|0.28|0.648|0.072|"RT @smoothkobra: A white Trump supporter just killed two cops and #BlueLivesMatter is nowhere to be found. They just hate Black people, tha"
fkatitle|hisillusion|0.5574|0.0|0.685|0.315|RT @hisillusion: Person: How does a typical Trump supporter look like? Me: https://t.co/sseV3ExOP5
fkatitle|twitter|0.5574|0.0|0.685|0.315|RT @hisillusion: Person: How does a typical Trump supporter look like? Me: https://t.co/sseV3ExOP5
CarlToddHand|jaynordlinger|0.4404|0.0|0.884|0.116|RT @jaynordlinger: If Bill Clinton talked Donald Trump into running for the GOP nomination -- Clinton truly is the wiliest politician in wo
yesbihjapril|Bill_Nye_Tho|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
yesbihjapril|twitter|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
clintonchineduc|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana 0.6% reporting TRUMP 69.8% | Hillary 26.4%  massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Elect
mxdelinneee|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
mxdelinneee|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
Brendag38323989|Sausage_House|0.5399|0.0|0.868|0.132|"RT @Sausage_House: Hey #Bernie supporters. Think about it. If you vote for Trump now, you'll only have to wait 4 years to try again!! https"
FehlJohn|TheLastRefuge2|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
FehlJohn|twitter|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
beltranaminta|HaskelBiz|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
beltranaminta|twitter|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
bea_nyce|Rivercasino7|-0.6059|0.205|0.728|0.068|"RT @Rivercasino7: Let me get this straight.. A MAN can punch, and throw a WOMAN down to the ground for supporting Trump, but no arrest is m"
Mongo10|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
stmpinfortrump|ilovemyfreedom|0.0|0.0|1.0|0.0|Rural Kentucky chimes in for TRUMP! https://t.co/3c1iOFyNSZ https://t.co/Wm05VnJkVe
revsaint08|drewwyatt|-0.5216|0.151|0.849|0.0|RT @drewwyatt: Hillary Campaign Paid Rioters 2 Burn The American Flag @ Trump Rally.You Can't Love Our Country &amp; Justify Voting 4 Her.
__sweetliar|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
__sweetliar|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
for_congress|AmericaFirst16|0.0|0.0|1.0|0.0|RT @AmericaFirst16: @FoxNews Votes are coming in KY and Ind and Trump is up FIFTY!Stop the BS #ElectionNight
beltranaminta|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
darcy027027|0hour|0.0|0.0|1.0|0.0|RT @0hour: Paris Hilton voted Trump BTFO!
gnoh_sandra|Jenn_Abrams|0.3612|0.0|0.783|0.217|RT @Jenn_Abrams: Donald Trump's web-site now looks like that https://t.co/s1yg0IthfJ
gnoh_sandra|twitter|0.3612|0.0|0.783|0.217|RT @Jenn_Abrams: Donald Trump's web-site now looks like that https://t.co/s1yg0IthfJ
56jaytee|costareports|0.4019|0.0|0.847|0.153|"RT @costareports: Kellyanne Conway to @chucktodd: Trump didnt have the full support of the Republican infrastructure"""
MarcusFromWV|.|0.0|0.0|1.0|0.0|If I was Trump I'd have entertainable people to Tweet @. Instead I have 154 followers who probably joined in 2008 &amp; forgot they have Twitter
tayleigh007|WDFx2EU8|0.8443|0.0|0.597|0.403|"RT @WDFx2EU8:  BREAKING: WOW!!! At the last minute, Chris Matthews endorses #Trump!!! #ElectionDay  https://t.co/FjeNWIsACt"
tayleigh007|twitter|0.8443|0.0|0.597|0.403|"RT @WDFx2EU8:  BREAKING: WOW!!! At the last minute, Chris Matthews endorses #Trump!!! #ElectionDay  https://t.co/FjeNWIsACt"
Down4Sue|jchesney266|0.4168|0.084|0.724|0.192|RT @jchesney266: @realDonaldTrump @jchesney266 @ScottPresler @mitchellvii Now this is a hard core Trump fan!!! https://t.co/SCeFNBVZab
Down4Sue|twitter|0.4168|0.084|0.724|0.192|RT @jchesney266: @realDonaldTrump @jchesney266 @ScottPresler @mitchellvii Now this is a hard core Trump fan!!! https://t.co/SCeFNBVZab
vmvanmoppes|GeorgeTakei|0.0|0.0|1.0|0.0|"RT @GeorgeTakei: Wait, wait. ""At least"" 4 grandparents? Just how many are we expected to have? We're not all Trump children with three poss"
inputfunction|jko417|0.0|0.0|1.0|0.0|"RT @jko417: ""Donald Trump is not the person that the media has depicted him to be"" #Trump2016 (Vine by @USAforTrump2016) https://t.co/R3G7K"
inputfunction|t|0.0|0.0|1.0|0.0|"RT @jko417: ""Donald Trump is not the person that the media has depicted him to be"" #Trump2016 (Vine by @USAforTrump2016) https://t.co/R3G7K"
Pfro|goldengateblond|-0.7184|0.222|0.778|0.0|RT @goldengateblond: The Trump campaign asked a judge to make the names of Nevada poll workers public. She had no time for their bullshit.
wtmkylie|brosemaiman|0.6486|0.0|0.739|0.261|@brosemaiman tomorrow @ school I have to debate with a trump supporter about health care &amp; I DONT WANNA GET ROASTED
kirtymom|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
kirtymom|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
littleicedragon|KeetPotato|0.5423|0.057|0.766|0.177|"RT @KeetPotato: [if trump wins somehow]alien: ""i said take me to your leader""me: ""dude i swear this is him"""
Woke_Silence|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
Woke_Silence|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
nothing_exists|chrislhayes|-0.5256|0.159|0.841|0.0|RT @chrislhayes: Trump is already laying the groundwork to contest the legitimacy of the election and it's incredibly dangerous.
This_is_ian_|SortaBad|-0.5423|0.132|0.868|0.0|"RT @SortaBad: Long line at this polling station, and it appears people are casting their votes in Spanish (soy, grande, etc). Bad sign for"
cr100064|WeNeedTrump|-0.5574|0.153|0.847|0.0|"RT @WeNeedTrump: By wanting to shut down illegal immigrantion, the Democrats and mainstream media have done everything possible to paint Tr"
deedemayo|Olivia_Baum|-0.7269|0.332|0.553|0.115|"RT @Olivia_Baum: If you support Trump, I consider you racist, sexist, and someone who condones sexual assault."
choozurlife|damaninthearena|0.0|0.0|1.0|0.0|RT @damaninthearena: @Vendetta92429 @antimarxis_ this map is BS!! I'm in southern Cali and in a line of 50+ people; Black White Hispanic As
Lane_bristow|gymstarz1053|-0.296|0.355|0.645|0.0|@gymstarz1053 no just vote trump
CarlosIsCarLost|MaduroOfficial|0.0|0.0|1.0|0.0|RT @MaduroOfficial: USA ELECTION UPDATEDonald Trump -   22.4%Hilary Clinton -   16.6%PSUV.               -  61.1%
xMOLONLABEx|hboulware|0.8555|0.0|0.606|0.394|"@hboulware Yes, I'm sure it was the same ""data"" sources that said Trump had a 1% chance of winning the primary...@ThomasPayne49"
lb_ashtoo|Kilerpollo78|-0.5423|0.28|0.72|0.0|RT @Kilerpollo78: Fuck Trump idc what any of yall say
KramerFry|nanodoug|0.5719|0.0|0.812|0.188|"RT @nanodoug: WIKILEAKS 1-35 BREAKING NEWS: Donald Trump Wins Florida, OH, NC Despite ... https://t.co/tYj4cJyKKH via @YouTube"
KramerFry|youtube|0.5719|0.0|0.812|0.188|"RT @nanodoug: WIKILEAKS 1-35 BREAKING NEWS: Donald Trump Wins Florida, OH, NC Despite ... https://t.co/tYj4cJyKKH via @YouTube"
givenchybey|rainymondays|0.0|0.0|1.0|0.0|RT @rainymondays: me to 'gays for trump' when i get sent to concentration camps &amp; see them there https://t.co/EI2nKmmPse
givenchybey|twitter|0.0|0.0|1.0|0.0|RT @rainymondays: me to 'gays for trump' when i get sent to concentration camps &amp; see them there https://t.co/EI2nKmmPse
ohmyswift1213|vibeeeez|-0.5574|0.261|0.739|0.0|RT @vibeeeez: prediction: Hillary Clinton is our next present &amp; everyone is shocked Trump lost
lexi_havel97|MaggieBecka|0.0258|0.113|0.769|0.117|RT @MaggieBecka: i am freaking the heck out over this election. i cannot understand why anyone would think trump would be a good leader
PsycGrrrl|Nebula63|0.4133|0.14|0.664|0.196|RT @Nebula63: Text to family: Don't expect me to be civil w any Trump supporters at any family gathering. Feel free to not invite me. I won
BaselGooner|larrymeath|-0.0276|0.093|0.818|0.089|RT @larrymeath: It's difficult to sneer at a nation who may very well put #Trump in White House   when your own nation has Boris Johnson a
tamaraleighllc|JoeyArnoldVN|0.0|0.0|1.0|0.0|RT @JoeyArnoldVN: GO VOTE TODAY TRUMP HILLARY CLINTON#ExitPoll#iVoted#myVote2016#ElectionDay#VoteJSA#Poll#WTFAmericaIn5Words#DolanT
TruthSmackdown|mitchellvii|0.4404|0.0|0.805|0.195|"RT @mitchellvii: Trump leads IND 72-25.  Good Lord people, something is happening here."
pattywc|cnnbrk|-0.4767|0.22|0.78|0.0|RT @cnnbrk: Eric Trump may have broken law with ballot tweet.  https://t.co/3cEkwFgO3p
pattywc|cnn|-0.4767|0.22|0.78|0.0|RT @cnnbrk: Eric Trump may have broken law with ballot tweet.  https://t.co/3cEkwFgO3p
_ayannnaaaa|ItsMeGrizz|-0.6124|0.154|0.846|0.0|RT @ItsMeGrizz: What is the real difference between Clinton and Trump for Black Ppl? Will either make steps to ending police brutality towa
taytay007007007|HalleyBorderCol|0.7703|0.0|0.74|0.26|"RT @HalleyBorderCol: For anyone wanting election results as them come in, the Guardian site seems quite good. Looking good for #Trump!htt"
Michaela_Govea|BlendlessBarlos|-0.8625|0.377|0.533|0.09|"RT @BlendlessBarlos: If you/ your parents support Donald trump fuck you , yo momma, yo grandmama &amp; fuck your dead homies"
iSoyJoel_|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
iSoyJoel_|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
junkyarddog66|reidepstein|0.6037|0.0|0.67|0.33|RT @reidepstein: A Trump runaway in Millsfield NH - 16-4 https://t.co/t1zLwKIhha
junkyarddog66|twitter|0.6037|0.0|0.67|0.33|RT @reidepstein: A Trump runaway in Millsfield NH - 16-4 https://t.co/t1zLwKIhha
valandspence|umpire43|0.2023|0.11|0.719|0.171|RT @umpire43: 2 Clinton supporters tried to bully me in line because of my Chemo hookup.Another Clinton supporter came to my aid then he vo
karenhunter|SXMUrbanView|0.0|0.0|1.0|0.0|RT @SXMUrbanView: History on Repeat: Trump Campaign Eerily Echoes Segregationist George Wallace https://t.co/NR5tiXPI9X @karenhunter Show #
karenhunter|atlantablackstar|0.0|0.0|1.0|0.0|RT @SXMUrbanView: History on Repeat: Trump Campaign Eerily Echoes Segregationist George Wallace https://t.co/NR5tiXPI9X @karenhunter Show #
Tehpanga|slayinglooks|0.0|0.0|1.0|0.0|RT @slayinglooks: Will Hillary make pants suits mandatory?Will Trump build a wall on Mexicos border?   Find out tomorrow on the season
webcentraltv|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
webcentraltv|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
IamtheCarmen__|Sportsmanshipp|0.0|0.0|1.0|0.0|RT @Sportsmanshipp: Gisele Refutes Donald Trump's Claim That Tom Brady Voted For Him https://t.co/0cF91sY8x4
IamtheCarmen__|12up|0.0|0.0|1.0|0.0|RT @Sportsmanshipp: Gisele Refutes Donald Trump's Claim That Tom Brady Voted For Him https://t.co/0cF91sY8x4
Roryyy_b|bet365|0.8225|0.0|0.703|0.297|Get trump to win the election at 9/2 or Clinton 1/6Underdog got the brexit win will it happen again? https://t.co/zvD2gTWU4I
redskinsrock91|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
ADrunkStitch|twitter|0.6449|0.0|0.652|0.348|Proud of mom for voting for Trump!!!!!! #FoxNews2016 https://t.co/u5hwNAssep
janna926|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump now leading IN by 45 points.  RCP has him by 10.  Something is happening.
DarrenRobyAZ|BlissTabitha|-0.4588|0.188|0.813|0.0|RT @BlissTabitha: Nevada Poll Workers Break Law: Caught Wearing Defeat Trump T-Shirts https://t.co/Ibt0aR0n4h #Election2016
DarrenRobyAZ|thegatewaypundit|-0.4588|0.188|0.813|0.0|RT @BlissTabitha: Nevada Poll Workers Break Law: Caught Wearing Defeat Trump T-Shirts https://t.co/Ibt0aR0n4h #Election2016
nct_doyoungg|greysonchance|-0.126|0.102|0.817|0.082|RT @greysonchance: To every American 18+...Go VOTE tomorrow! We have a chance to stop Donald Trump from ever stepping into the Oval Office
dejean76|gerfingerpoken|0.0|0.0|1.0|0.0|"RT @gerfingerpoken: Trump Defends Life, Hillary Defends #PartialBirthAbortion - Flopping Aces - https://t.co/boHSpqQIqN #MAGA https://t.co/"
dejean76|floppingaces|0.0|0.0|1.0|0.0|"RT @gerfingerpoken: Trump Defends Life, Hillary Defends #PartialBirthAbortion - Flopping Aces - https://t.co/boHSpqQIqN #MAGA https://t.co/"
vision835|twitter|0.0|0.0|1.0|0.0|TRUMP! https://t.co/nH9DG6nxbW
peaceoutanddab|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
crose84|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
crose84|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
SupaKawaiiLexi|ScienceTrash|0.4201|0.0|0.877|0.123|"@ScienceTrash But it still has to go through Congress. I'm not for Trump, or Hillary. So I agree with what you're saying."
donna_heinrich|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
__hamishh|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
forphiI|chokemehowelI|-0.4023|0.172|0.828|0.0|RT @chokemehowelI: rt this if you wouldnt feel comfortable sitting in a room with trump
VilleSZN|JayeNick_|-0.5719|0.236|0.764|0.0|RT @JayeNick_: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/dpWCWHwHhw
VilleSZN|twitter|-0.5719|0.236|0.764|0.0|RT @JayeNick_: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/dpWCWHwHhw
HopeSlick|JamilahLemieux|-0.2732|0.087|0.87|0.043|"RT @JamilahLemieux: No matter what happens tonight, the fact that Donald Trump has gotten this far is a stain on America that can't be wash"
DNoticie|ilovemyfreedom|0.0|0.0|1.0|0.0|Rural Kentucky chimes in for TRUMP! https://t.co/BH2oyRWM7S https://t.co/17mx8copIt
societygirl123|2ALAW|0.0|0.0|1.0|0.0|RT @2ALAW: Donald Trump #FoxNews2016 #electionday https://t.co/SI37Q8hESv
societygirl123|twitter|0.0|0.0|1.0|0.0|RT @2ALAW: Donald Trump #FoxNews2016 #electionday https://t.co/SI37Q8hESv
CKlein5852|AdamsFlaFan|-0.128|0.215|0.633|0.152|RT @AdamsFlaFan: Hero Judge Stands Up For Democracy And Rejects Trump's Nevada Election Day Lawsuit via @politicususa https://t.co/v32RI9gi
CKlein5852|t|-0.128|0.215|0.633|0.152|RT @AdamsFlaFan: Hero Judge Stands Up For Democracy And Rejects Trump's Nevada Election Day Lawsuit via @politicususa https://t.co/v32RI9gi
brandvoldemort|DeanteVH|0.0|0.0|1.0|0.0|RT @DeanteVH: Trump can't run his own Twitter but people think he can run a country. Y'all wild https://t.co/5xZPUykUyJ
brandvoldemort|twitter|0.0|0.0|1.0|0.0|RT @DeanteVH: Trump can't run his own Twitter but people think he can run a country. Y'all wild https://t.co/5xZPUykUyJ
R_Kirun1|Fusion|-0.128|0.113|0.795|0.092|"RT @Fusion: ""Since he's gonna lose, I'm going to go dancing.""Latinas share #ElectionNight predictions at the Nevada store Trump tried &amp; f"
laurajeannee|chlolowin|0.0|0.0|1.0|0.0|RT @chlolowin: Why would anyone in their right mind vote for Donald Trump??? #ElectionDay
UwuaMan|RollingStone|0.34|0.0|0.87|0.13|"See Bruce Springsteen Play Solo, Rip Trump at Clinton Rally https://t.co/nyS4Dgnc7u via @RollingStone #uwua #labor #union #unions"
UwuaMan|rollingstone|0.34|0.0|0.87|0.13|"See Bruce Springsteen Play Solo, Rip Trump at Clinton Rally https://t.co/nyS4Dgnc7u via @RollingStone #uwua #labor #union #unions"
Dreamchasers_15|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Dreamchasers_15|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
sluggoD54|peaceandjoy101|0.6908|0.0|0.787|0.213|RT @peaceandjoy101: By asking Durham County North Carolina voting polls to remain open until 9pm is a sure sign Trump is winning in NC.#El
LeahR77|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
junebugjeanne|LynnKuennen|0.8225|0.0|0.743|0.257|RT @LynnKuennen: BREAKING: Trump on Hannity:  If we get panhandle and I40 corridor out to vote tonight we win Florida.  We can win Michigan
mstazrn|kachninja|0.0|0.0|1.0|0.0|"RT @kachninja: Just voted!!! #MAGA3X  My MIL went with us, a reformed Democrat for Trump!!! #IVotedTrump #VotingDay https://t.co/55oZJkYH"
mstazrn|t|0.0|0.0|1.0|0.0|"RT @kachninja: Just voted!!! #MAGA3X  My MIL went with us, a reformed Democrat for Trump!!! #IVotedTrump #VotingDay https://t.co/55oZJkYH"
blkshirtfan|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
kaylaabarness|BernieSanders|0.4404|0.113|0.68|0.207|RT @BernieSanders: Donald Trump is proud of his assaults on women and makes fun of people with disabilities. That is not someone who should
jmeclk|LEFTH00K|0.0|0.0|1.0|0.0|"RT @LEFTH00K: BREAKING: For the first time EVER more than 40,000 AMISH in PENNSYLVANIA will VOTE &amp; VOTE FOR TRUMP!20 BUSES TAKING THEM TO P"
sulamifschukin5|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
sulamifschukin5|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
CaldoHendo|rblandford|-0.5574|0.31|0.69|0.0|RT @rblandford: Shit. Sunderland South have gone for Trump.
CarolinaKT|THETXEMBASSY|0.0|0.0|1.0|0.0|@THETXEMBASSY #Trump will be our 45th President
InfamousVirgo|AriBerman|0.4404|0.0|0.873|0.127|RT @AriBerman: UPDATE: police came to polling place &amp; got control of situation. Trump supporters now off to the side https://t.co/bgn489aKsp
InfamousVirgo|twitter|0.4404|0.0|0.873|0.127|RT @AriBerman: UPDATE: police came to polling place &amp; got control of situation. Trump supporters now off to the side https://t.co/bgn489aKsp
iIoveharry|yvezayntIaurent|-0.5423|0.22|0.78|0.0|"RT @yvezayntIaurent: white person: idk whos worse: hillary or trumplgbtq, women, black people, immigrants, muslims: trump iswhite pers"
jewelagave|Hisladydiana|0.6114|0.0|0.693|0.307|RT @Hisladydiana: #Trump Our new President. America loves you ! https://t.co/l3Ix0dyxrx
jewelagave|twitter|0.6114|0.0|0.693|0.307|RT @Hisladydiana: #Trump Our new President. America loves you ! https://t.co/l3Ix0dyxrx
bryceMartian54|memetribute|-0.1695|0.186|0.814|0.0|"RT @memetribute: We don't want Trump, we don't want Hillary, we just want Cory back in the house #ElectionDay"
DaviGont|ESPACOAGRESSIVO|-0.6408|0.514|0.486|0.0|RT @ESPACOAGRESSIVO: FUCK TRUMP. https://t.co/VBIWEiQfYX
DaviGont|twitter|-0.6408|0.514|0.486|0.0|RT @ESPACOAGRESSIVO: FUCK TRUMP. https://t.co/VBIWEiQfYX
JDE6321|iResistAll|0.6249|0.0|0.779|0.221|"RT @iResistAll: BREAKING: Durham County, NC to extend voting in Democrat areas because Trump is winning the state. #electionday #ElectionN"
trapgod349|LouieVRee|-0.8271|0.3|0.636|0.064|RT @LouieVRee: Trump gay as hell if he trying to get rid of all the fine big booty Latina bitches too
annaklineee15|jessikab72|-0.5719|0.171|0.829|0.0|"RT @jessikab72: Remember: Trump has Pence, and he's enough of a reason to vote trump even if you hate trump"
samrobinson_96|mistry223|0.0|0.0|1.0|0.0|RT @mistry223: If the UK leaves the EU and Trump becomes president of the US in the same year I'm going to India to farm cows and make chee
marideenow|SimretZeru|0.0|0.0|1.0|0.0|"RT @SimretZeru: ""@MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/G9IQjfWImd"" #Canada"
marideenow|twitter|0.0|0.0|1.0|0.0|"RT @SimretZeru: ""@MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/G9IQjfWImd"" #Canada"
Brain1Brain|BiancaJagger|-0.6369|0.279|0.615|0.107|"RT @BiancaJagger: Dear Jon Donald Trump is not only a sociopath, he is a racist, xenophobic and a women hater https://t.co/E6D1i3aSPr"
Brain1Brain|twitter|-0.6369|0.279|0.615|0.107|"RT @BiancaJagger: Dear Jon Donald Trump is not only a sociopath, he is a racist, xenophobic and a women hater https://t.co/E6D1i3aSPr"
_kyanaaaa|twitter|0.5106|0.0|0.476|0.524|Free Teanna Trump  https://t.co/RkGhFmmlpR
ReaganBattalion|twitter|0.7184|0.0|0.4|0.6|Still 100% sure Trump wins? https://t.co/AYkFaMoIVZ
BoycottHRC|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
pandaonparole|CNN|0.3182|0.0|0.881|0.119|@CNN even when he dies the DemocRATS will make sure he still casts his vote #VoterFraud #Trump #MakeAmericaGreatAgain
LeoReynaJr|jpodhoretz|-0.1531|0.091|0.909|0.0|"RT @jpodhoretz: Sara Murray on CNN says Trump source says a ""key internal metric"" shows Trump falling short"
negative_niko|fivethirtyeight|0.2023|0.196|0.515|0.289|Good article about bullshit narrative of Trump's support being majority working class https://t.co/OB4ehekE4c
party_poisonous|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
party_poisonous|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
iSydneyNews|christianitytoday|0.2023|0.0|0.886|0.114|Top 10 Stats Explaining the Evangelical Vote for Trump or Clinton https://t.co/Geo3lHIwMC #Sydney #News #Aus
twdmaIum|ObamaSpotify|-0.5423|0.226|0.774|0.0|RT @ObamaSpotify: President Obama is currently listening to Fuck Donald Trump by YG
jamiegirl|pewdrdad|0.4404|0.0|0.847|0.153|"RT @pewdrdad: First Early Exit Polls Just Released, and They Point Towards Good News for Trump https://t.co/ecsrFIRiXj"
jamiegirl|pinterest|0.4404|0.0|0.847|0.153|"RT @pewdrdad: First Early Exit Polls Just Released, and They Point Towards Good News for Trump https://t.co/ecsrFIRiXj"
cissysphotos|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
SportsInsights|twitter|0.0|0.0|1.0|0.0|Current #Florida Odds (Bookmaker)Clinton -319Trump +266#ElectionNight https://t.co/DVEtfn7nkK
Zoom81|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
thadarktruth|mcuban|0.0243|0.11|0.776|0.114|@mcuban I like how you offered Trump 10million to explain his policies and he didn't take the easy money. SMH...
NancyNielsenn|marwilliamson|0.0|0.0|1.0|0.0|@marwilliamson GO Trump!
SheenaMarie412|GeorgeTakei|0.0|0.0|1.0|0.0|"RT @GeorgeTakei: Of course, this would also disqualify Trump himself, whose grandparents were ALL born outside the USA... https://t.co/IIZs"
SheenaMarie412|t|0.0|0.0|1.0|0.0|"RT @GeorgeTakei: Of course, this would also disqualify Trump himself, whose grandparents were ALL born outside the USA... https://t.co/IIZs"
TrumpWithUSA|NeilTurner_|0.0516|0.125|0.741|0.134|RT @NeilTurner_: #VoterFraud Funny how there never seems to be issues with choosing #CrookedHillary. Always problems choosing Trump.#El
joannele2001|LadyLibertyWDC|0.0|0.0|1.0|0.0|RT @LadyLibertyWDC: Kentucky's got it going for Trump! https://t.co/Q8gA7KOcEG
joannele2001|twitter|0.0|0.0|1.0|0.0|RT @LadyLibertyWDC: Kentucky's got it going for Trump! https://t.co/Q8gA7KOcEG
Make_Me_Smil3|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Make_Me_Smil3|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
notericisboss84|BoofBaldy|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
notericisboss84|twitter|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
Hanto38Le|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
Hanto38Le|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
KristinaF1977|FreddieCampion|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
KristinaF1977|twitter|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
Megmo808|ErickFernandez|-0.4019|0.171|0.829|0.0|RT @ErickFernandez: Nevada judge did not have time for Trump's lawsuit complaining that too many brown people voted. #ElectionDay https://t
Megmo808||-0.4019|0.171|0.829|0.0|RT @ErickFernandez: Nevada judge did not have time for Trump's lawsuit complaining that too many brown people voted. #ElectionDay https://t
SmitaRanjit|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
SmitaRanjit|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
RoniSeale|joelpollak|0.4019|0.0|0.838|0.162|RT @joelpollak: Trump Fans Sing Star-Spangled Banner in Front of Victory Party https://t.co/wVlNFT9hzp via @BreitbartNews
RoniSeale|breitbart|0.4019|0.0|0.838|0.162|RT @joelpollak: Trump Fans Sing Star-Spangled Banner in Front of Victory Party https://t.co/wVlNFT9hzp via @BreitbartNews
Life_Force_1|twitter|0.0|0.0|1.0|0.0|REPEAT AFTER ME:  DONDALD J TRUMP WILL BE PRESIDENT #Decision2016 #MAGA3X #GlobalShift #TRUMP https://t.co/V8OQSEekIg
Aspennicole17|precious_oxox|-0.6169|0.314|0.686|0.0|RT @precious_oxox: this election is fucking with my anxiety. Donald Trump cannot win.
pablo_pachecoo|FableofJosh|-0.1027|0.149|0.851|0.0|RT @FableofJosh: Trump: *loses*Trump: nah I never ran for president
ramesh_tnt|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
ramesh_tnt|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
Axellent33|Verge|0.5106|0.0|0.708|0.292|Donald Trump's website enjoyed a brief democracy https://t.co/y7zBMbqU8i via @Verge
Axellent33|theverge|0.5106|0.0|0.708|0.292|Donald Trump's website enjoyed a brief democracy https://t.co/y7zBMbqU8i via @Verge
endeeh|speechboy71|-0.5106|0.202|0.798|0.0|RT @speechboy71: If only Trump had insulted the spouses of every Republican #whatcouldhavebeen https://t.co/ElY8QxJL3U
endeeh|twitter|-0.5106|0.202|0.798|0.0|RT @speechboy71: If only Trump had insulted the spouses of every Republican #whatcouldhavebeen https://t.co/ElY8QxJL3U
Angelmdunn1961|Democrat_4Trump|0.6249|0.0|0.819|0.181|RT @Democrat_4Trump: Poll closing by STATE.Get out and vote if you haven't done so yet. Trump NEEDS EVERY VOTE. We want to win folks. @rea
bavcena66|CJMatthews25|0.7177|0.0|0.778|0.222|Hey @CJMatthews25 can you warm up a bed in case Trump manages to win? I already know the Canadian national anthem in English &amp; French!
JimJesus|youtube|0.4019|0.0|0.803|0.197|Tonight we watch Trump burn the Republican Party to the ground. https://t.co/CQQizBGR3X
killahectaa|rainymondays|0.0|0.0|1.0|0.0|RT @rainymondays: me to 'gays for trump' when i get sent to concentration camps &amp; see them there https://t.co/EI2nKmmPse
killahectaa|twitter|0.0|0.0|1.0|0.0|RT @rainymondays: me to 'gays for trump' when i get sent to concentration camps &amp; see them there https://t.co/EI2nKmmPse
MishaMishaps|kurteichenwald|-0.4033|0.244|0.609|0.147|"RT @kurteichenwald: I just realized: With Nevada, Trump is essentially arguing that allowing people to vote is voter fraud. Quite amazing w"
Matiias_Denmon|smoothkobra|-0.7964|0.28|0.648|0.072|"RT @smoothkobra: A white Trump supporter just killed two cops and #BlueLivesMatter is nowhere to be found. They just hate Black people, tha"
erik_dvoxo|gar_gar21|0.25|0.0|0.882|0.118|RT @gar_gar21: I had a dream I voted for Donald Trump last night.. scariest nightmare I've had in months
ItsThatGuyBrent|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
ItsThatGuyBrent|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
MsHoefler|chrislhayes|0.0|0.0|1.0|0.0|"RT @chrislhayes: After waiting until almost *literally* the last moment, Toomey votes and says he voted for Trump."
JulieCTaylor|twitter|0.5859|0.0|0.833|0.167|Amazing that I never see reports of votes switching from Hillary to Trump. Always the other way. Makes me wonder.Hm https://t.co/yu85qCqIYp
sanchez03h|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
sanchez03h|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
citroncool|dril|0.0|0.0|1.0|0.0|RT @dril: if you ask me this election could end about 100 different ways:1) trump gets 0% of the vote2) trump gets 1% of the vote3) trum
marveItrade|mashable|0.0|0.0|1.0|0.0|RT @mashable: Caught! Donald Trump was peeking at his wife's election ballot  #ElectionNight https://t.co/1CsOJNnkpo
marveItrade|twitter|0.0|0.0|1.0|0.0|RT @mashable: Caught! Donald Trump was peeking at his wife's election ballot  #ElectionNight https://t.co/1CsOJNnkpo
joehanraty|BlueyezEST|0.0|0.0|1.0|0.0|"RT @BlueyezEST: TWITTER POLL, WHO WILL BE THE NEXT U.S PRESIDENT? #trump #clinton #ElectionDay #ElectionNight #PresidentialElection2016 #Do"
trading24h|RampCapitalLLC|0.34|0.0|0.854|0.146|RT @RampCapitalLLC: Excited for a MSM meltdown if Trump carries a lead for more than an hour
franklapore|politico|-0.5859|0.348|0.652|0.0|Trump seizes on isolated glitches to fuel rigged election claims  https://t.co/AVEY0b9tPT
FedoraPayan|NicoleG5555|0.25|0.117|0.676|0.207|RT @NicoleG5555: @bea_nyce @wesearchr @reddit @FoxNews @foxandfriends Trump will fight This. Thank God for the videos.  #riggedelection #Ri
Stepto|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
EricStoller|thenation|0.0|0.0|1.0|0.0|Dont Tell Trump: Minnesota Is About to Elect a Pioneering Somali-American Muslim Woman | #Election2016  https://t.co/tgmKtrHXA7
CortocircuitOFi|mazthetelling|0.6249|0.0|0.745|0.255|RT @mazthetelling: Great - Hop Frog FB: https://t.co/6BWcAPaU9n #ElectionDay #ElectionNight #Trump #maratonamentana @DinamoPress https://t.
CortocircuitOFi|m|0.6249|0.0|0.745|0.255|RT @mazthetelling: Great - Hop Frog FB: https://t.co/6BWcAPaU9n #ElectionDay #ElectionNight #Trump #maratonamentana @DinamoPress https://t.
Nandobyson28|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
Cavalli512|VAWSE|0.0|0.0|1.0|0.0|RT @VAWSE: YESSSS RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/JuZm7ayVoY
Cavalli512|twitter|0.0|0.0|1.0|0.0|RT @VAWSE: YESSSS RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/JuZm7ayVoY
tomseward|peddoc63|0.3182|0.0|0.905|0.095|"RT @peddoc63: My 19 year old son 1st supported Bernie Sanders, then Gary Johnson, today he is voting for Donald J. Trump#ElectionNight #m"
Alinglese|JimSavell|0.0|0.0|1.0|0.0|RT @JimSavell: @catoletters Have you seen the videos of people not being able to vote for Trump? They click the button and nothing happens
BrendaGL9|DaniellBautista|-0.6408|0.458|0.542|0.0|RT @DaniellBautista: FUCK DONALD TRUMP https://t.co/0TUaRyRjgJ
BrendaGL9|twitter|-0.6408|0.458|0.542|0.0|RT @DaniellBautista: FUCK DONALD TRUMP https://t.co/0TUaRyRjgJ
neyotherock|TrustedKenyan|-0.4023|0.153|0.847|0.0|RT @TrustedKenyan: Donald Trump doesn't trust his wife Maybe he dreamt her voting for Clinton https://t.co/7bbjV0FRvA
neyotherock|twitter|-0.4023|0.153|0.847|0.0|RT @TrustedKenyan: Donald Trump doesn't trust his wife Maybe he dreamt her voting for Clinton https://t.co/7bbjV0FRvA
wondaland|BetteMidler)I|-0.5852|0.226|0.774|0.0|Retweeted Bette Midler (@BetteMidler):I guess the Trump men don't really trust their wives!!!... https://t.co/BNOFfDyIur
wondaland|twitter|-0.5852|0.226|0.774|0.0|Retweeted Bette Midler (@BetteMidler):I guess the Trump men don't really trust their wives!!!... https://t.co/BNOFfDyIur
PatsSoxBruins|C_Danielle16|-0.567|0.197|0.803|0.0|@C_Danielle16 trump then I am sorry you have participated in not wanting to preserve our planet for future generations  Just so upset
SynergyByDesign|EmilyMiller|0.4574|0.0|0.857|0.143|RT @EmilyMiller: I'll be live on @OANN all #ElectionNight from Trump NYC party. Tune in for the latest! https://t.co/umIpjVDrjO
SynergyByDesign|twitter|0.4574|0.0|0.857|0.143|RT @EmilyMiller: I'll be live on @OANN all #ElectionNight from Trump NYC party. Tune in for the latest! https://t.co/umIpjVDrjO
ttm2x|DJ_SKEME|0.7579|0.0|0.629|0.371|RT @DJ_SKEME: #BlackTwitter will be pure entertainment tonight whether Hillary or Trump wins
Beachbored2|mr_kyloving|-0.2263|0.142|0.751|0.107|"RT @mr_kyloving: Rob O Neil ""98% of U.S special forces are voting Trump"" the other 2% are going for Gary Johnson. @realDonaldTrump"
knew777771|LOLGOP|0.0516|0.138|0.714|0.148|RT @LOLGOP: EXIT POLL: 3 in 10 Trump supporters had trouble finding the exit to the polls.
MayorSnart|Queentette|0.5996|0.069|0.701|0.23|@Queentette Hillary isn't a white straight male. So everything she does is ok. As long as she's not that scumbag Trump
amuses|DonaldJTrumpJr|0.8398|0.0|0.69|0.31|"RT @DonaldJTrumpJr: Please watch and share this. Vote now to take back America! ""Freedom is never more than one generation away from exti"
getalifegoldy|Teckerke|-0.5439|0.392|0.608|0.0|@Teckerke probably some crazy person how didnt like trump
Ddubb__|HillaryClinton|0.2382|0.143|0.64|0.217|I don't give a fuck about none of these Trump supporters cause regardless my bitch @HillaryClinton finna come out with this dub
NJHomesKOOLMom|davidplouffe|0.4404|0.0|0.756|0.244|@davidplouffe @JanetMenke Your bar looks better than Trump's cash bar
ExitsRevolution|sciam|-0.2006|0.121|0.879|0.0|RT @sciam: Here are some of Donald Trump's most alarming statements about science https://t.co/Q4fD0zoPzw
ExitsRevolution|scientificamerican|-0.2006|0.121|0.879|0.0|RT @sciam: Here are some of Donald Trump's most alarming statements about science https://t.co/Q4fD0zoPzw
ARMY_PARENT|Thomas1774Paine|0.0|0.0|1.0|0.0|RT @Thomas1774Paine: Female #Trump voter hammers CNN. Yinz shouldn't have asked the question if Yinz at CNN didn't know the answer. Google
clutchdom23|twitter|0.0|0.0|1.0|0.0|"""You voting for Trump"" https://t.co/80Yo2x63dP"
216JDoeYahhh|YoungDems4Trump|-0.582|0.334|0.444|0.222|"@YoungDems4Trump I know for sure Trump supporters are angry Bernie didn't win because even if Trump lost, at least it was a fair fight."
KingPlaysClaw|ImPeacefulChaos|0.0|0.0|1.0|0.0|RT @ImPeacefulChaos: RT for this rockLike for Trump https://t.co/CvbTA8llrP
KingPlaysClaw|twitter|0.0|0.0|1.0|0.0|RT @ImPeacefulChaos: RT for this rockLike for Trump https://t.co/CvbTA8llrP
Linda_2008|LarrySchweikart|0.0|0.0|1.0|0.0|@LarrySchweikart trump jr was just on Hannity saying panhandle needs to go vote? Where did u get those #s
Amirez_CHARMS|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
Amirez_CHARMS|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
Koxinga8|breitbart|0.5859|0.0|0.774|0.226|Frank Luntz: #Trump Could Win Michigan  Working-Class Turnout 'Much Higher than Expected' - Breitbart https://t.co/gIclIzCOzS
ia_yeah|aidan|0.765|0.0|0.732|0.268|RT @aidan: trump showing up to his polling place and getting booed is honestly the funniest thing i've ever seen
EEGRC98|0hour|0.0|0.0|1.0|0.0|RT @0hour: Kentucky Trump 69% Lads!
wildwalkerwoman|KTEwing901|-0.2411|0.079|0.921|0.0|RT @KTEwing901: #ElectionDay Reminder: Black people are not responsible for the rise of Trump. We did not place him in this position. He is
sophia7213|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
jeanne_tall|Mike_Beacham|0.0|0.0|1.0|0.0|RT @Mike_Beacham: Donald Trump: The Candidate Who Never Quit @realDonaldTrump @DonaldJTrumpJr @EricTrump @IvankaTrump #MAGA #tcothttp
POPPER722|twitter|0.54|0.0|0.858|0.142|He's going to have plenty of time to talk to himself with his very good brain in solitary confinement! Trump Univer https://t.co/CX0LzEqjZk
davedbody|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
davedbody|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
kylesnooze|cracked|-0.0258|0.046|0.954|0.0|"RT @cracked: ""I've long awaited this,"" murmured Trump Jr., as he took a chunk of his father's cake face in his fist and squeeeezed. https:/"
kylesnooze||-0.0258|0.046|0.954|0.0|"RT @cracked: ""I've long awaited this,"" murmured Trump Jr., as he took a chunk of his father's cake face in his fist and squeeeezed. https:/"
paigeatzemis|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
paigeatzemis|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
cevenwebb76|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
cevenwebb76|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
tallysimone|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
tallysimone|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
VirgPatriot|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump now leading IN by 45 points.  RCP has him by 10.  Something is happening.
_lulshawtyyy|stayguccisam|0.6739|0.058|0.74|0.203|RT @stayguccisam: The hispanics voting for trump probably LOVE to pretend to be white and only speak English at home
Da1nOnlyCMart|KTLA|0.2732|0.0|0.89|0.11|"RT @KTLA: Clinton and Trump supporter exchange blows, pepper spray during scuffle at Florida polling site https://t.co/yRWvop7e1b https://t"
Da1nOnlyCMart|ktla|0.2732|0.0|0.89|0.11|"RT @KTLA: Clinton and Trump supporter exchange blows, pepper spray during scuffle at Florida polling site https://t.co/yRWvop7e1b https://t"
lilulyvert_|SOMEXlCAN|-0.4404|0.25|0.595|0.155|RT @SOMEXlCAN: YOOO SOMEONE PLAYED MEXICAN MUSIC AT A DONALD TRUMP RALLY IM DEAD  https://t.co/OJ2RJgfILk
lilulyvert_|twitter|-0.4404|0.25|0.595|0.155|RT @SOMEXlCAN: YOOO SOMEONE PLAYED MEXICAN MUSIC AT A DONALD TRUMP RALLY IM DEAD  https://t.co/OJ2RJgfILk
Sva98_|TakeSimplAdvice|0.5719|0.0|0.654|0.346|RT @TakeSimplAdvice: Trump voters if Trump wins https://t.co/YyvI4JHwxN
Sva98_|twitter|0.5719|0.0|0.654|0.346|RT @TakeSimplAdvice: Trump voters if Trump wins https://t.co/YyvI4JHwxN
DaddyMalena|jaketapper|0.3566|0.0|0.894|0.106|"RT @jaketapper: But then Trump couldn't run, since his mom and paternal grandparents weren't born in the US. So, um, yeah. https://t.co/7Ux"
DaddyMalena|t|0.3566|0.0|0.894|0.106|"RT @jaketapper: But then Trump couldn't run, since his mom and paternal grandparents weren't born in the US. So, um, yeah. https://t.co/7Ux"
ttsdunn|nationdivided|0.0|0.0|1.0|0.0|RT @nationdivided: Breaking news: @CNN is reporting that black turnout in Detroit is down 50% over 4 years ago that is Trump's pathway to w
theonlynoe|quuay__|0.0|0.0|1.0|0.0|"RT @quuay__: Only reason why white people voting for trump they think it's going to be how it was back in the days but,i think tf not."
chimmychann|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
chimmychann|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
BULGEBULL|i2|0.4019|0.0|0.838|0.162|WATCH LIVE: Hillary Clinton and Donald Trump Hold Election Night Parties Only A Mile Apart  https://t.co/vGY5zOkGg6
viplive|tmz|0.0|0.0|1.0|0.0|Hillary and Donald -- Enough Already!!! You're Bleeding Us Dry https://t.co/5pXLd0oILP
jmnphx|ShannonBream|0.5563|0.122|0.63|0.248|"@ShannonBream You fail to mention, the majority of trending ""Clinton"" on Facebook is negative.. While Trump is positive. You're very pretty."
Carolan2016|FoxNews|0.8159|0.0|0.547|0.453|@FoxNews RUSSIA READY FOR CLINTON PRESIDENCY   VOTE PEACE VOTE TRUMP  https://t.co/BUnS7SXwkJ
Carolan2016|rt|0.8159|0.0|0.547|0.453|@FoxNews RUSSIA READY FOR CLINTON PRESIDENCY   VOTE PEACE VOTE TRUMP  https://t.co/BUnS7SXwkJ
LabourNHSJAN|independent|0.296|0.0|0.885|0.115|Eric Trump illegally shares photo of him voting for his dad to be president | The Independent - www.independent. https://t.co/oee14c9qiI
bjw2112|mitchellvii|0.4648|0.0|0.664|0.336|"RT @mitchellvii: Again, HUGE FOR TRUMP. https://t.co/osXpZyBcze"
bjw2112|twitter|0.4648|0.0|0.664|0.336|"RT @mitchellvii: Again, HUGE FOR TRUMP. https://t.co/osXpZyBcze"
karbob85|hardassettimes|0.5719|0.0|0.793|0.207|RT @hardassettimes: @BarbMuenchen @maggiebeauchamp All those people are certainly not waiting in line to vote for Crooked Hillary. Pray for
OdellSZN|StephForMVP30|0.7955|0.0|0.718|0.282|RT @StephForMVP30: If Trump or Hillary wins the election I'm moving out the country! Goodbye America and hello United States!
garza16lisa|Bdell1014|0.0|0.0|1.0|0.0|RT @Bdell1014: I cant believe ppl are going to vote for a 70 year old man named Trump who had his twitter taken away cause he couldn't be t
smp0711|mtracey|0.0|0.0|1.0|0.0|"RT @mtracey: Former Sanders delegate from PA sends over this photo: voted Trump, then Democrats down ballot https://t.co/qfwbyhwIFx"
smp0711|twitter|0.0|0.0|1.0|0.0|"RT @mtracey: Former Sanders delegate from PA sends over this photo: voted Trump, then Democrats down ballot https://t.co/qfwbyhwIFx"
TylerHu99890202|FrankLuntz|0.25|0.0|0.889|0.111|RT @FrankLuntz: BREAKING: Watch Michigan.Working-class turnout is looking much higher than expected. Trump may actually have a chance.  #
seamusdf|ignitingflames|0.3885|0.157|0.581|0.262|"RT @ignitingflames: IDGI HOW ARE THERE PPL THAT SAY ""YEAH I DONT LIKE EITHER CANDIDATE BUT TRUMP IS BY FAR THE BETTER CANDIDATE"" YALL SCARY"
Doory25911|Democrat_4Trump|0.7269|0.0|0.711|0.289|RT @Democrat_4Trump: Current reporting in Kentucky and Indiana indicates a huge win for Trump. WATCH FOR #VoterFraud https://t.co/PWuqR6mmhS
Doory25911|twitter|0.7269|0.0|0.711|0.289|RT @Democrat_4Trump: Current reporting in Kentucky and Indiana indicates a huge win for Trump. WATCH FOR #VoterFraud https://t.co/PWuqR6mmhS
Wjk1027|HiHoblue22P|0.5411|0.0|0.845|0.155|RT @HiHoblue22P: #FrankLuntz did you notice how your Hand Picked Groups always get it Wrong!This Clinched IT for #Trump#TrumpTrain https:
Revitte||0.5267|0.0|0.694|0.306|"What #Trump &amp; his supporters are feeling now... @ Brooklyn, New York https://t.co/kM22JRBEPe"
Revitte|instagram|0.5267|0.0|0.694|0.306|"What #Trump &amp; his supporters are feeling now... @ Brooklyn, New York https://t.co/kM22JRBEPe"
sokolowski_g|realDonaldTrump|0.0|0.0|1.0|0.0|@realDonaldTrump @DonaldJTrumpJr I voted Trump!
laurie6805|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
laurie6805|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
Emylie|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
Emylie|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
backwaterdogs|mitchellvii|0.4404|0.0|0.838|0.162|"RT @mitchellvii: If Trump ends up dramatically outperfroming his RCP averages in early states, good sign."
PastorTeeTalley|wiselatinaslink|0.4019|0.0|0.863|0.137|RT @wiselatinaslink: Hillary Clinton will treat women as equals. You know what Trump thinks of us. #ElectionNight https://t.co/jgMQt6sGbk
PastorTeeTalley|twitter|0.4019|0.0|0.863|0.137|RT @wiselatinaslink: Hillary Clinton will treat women as equals. You know what Trump thinks of us. #ElectionNight https://t.co/jgMQt6sGbk
KweschnMedia|ajplus|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
KweschnMedia|twitter|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
EnidTheFairy|UnitatoCreation|0.5719|0.0|0.73|0.27|"RT @UnitatoCreation: If Trump wins, I'll draw everyone who rts this."
OccupyRadio3|news|0.0|0.0|1.0|0.0|How The Rest Of The World Sees Donald Trump: 12 Foreign Political Cartoons https://t.co/39FJc6VWth
AliceCoven|tommygunn12us|0.4404|0.0|0.674|0.326|RT @tommygunn12us: Looking good for trump. https://t.co/AqGBOVcG9X
AliceCoven|twitter|0.4404|0.0|0.674|0.326|RT @tommygunn12us: Looking good for trump. https://t.co/AqGBOVcG9X
Fullerforyotes|JoshuaCaudill85|-0.296|0.128|0.872|0.0|@JoshuaCaudill85 Syrian refugees are being properly vetted. Stop listening to trump. It's an extensive vetting system.
AliceCoven|ChooseToBFree|-0.7506|0.39|0.61|0.0|"RT @ChooseToBFree: @ezinder Aiding and abetting the enemy IS treason, Sir. @HlLLARYCLINT0N#HillaryIndictment#HillarysEmails#Hillary#Dra"
ChrisM_SF|benutty|-0.2235|0.173|0.827|0.0|"@benutty Trump's has a cash bar. Literally, that's not even a joke."
myidolismiranda|1432721|0.7626|0.0|0.477|0.523|@1432721 BECAUSE I DONT WANT TRUMP TO WIN THIS 
AriannaToledo23|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
AriannaToledo23|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Marcinzi|KevinGeb|0.4019|0.0|0.748|0.252|My Trump 2016 party about to be popping @KevinGeb
gia_mccomb|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
gia_mccomb|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
sassrin6|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
sassrin6|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
phenomenoire|surprise_bees|-0.4404|0.142|0.777|0.081|"RT @surprise_bees: It's like if Trump and Don Knotts fucked a cake, and that cake had a baby that grew old before its time and had seen too"
Redheadedbird|DiamondandSilk|0.3612|0.0|0.902|0.098|"RT @DiamondandSilk: If you are ready for Crooked Hill to EXIT then it's time for the American people to do a BREXIT.  ""Vote Trump"" https://"
Redheadedbird||0.3612|0.0|0.902|0.098|"RT @DiamondandSilk: If you are ready for Crooked Hill to EXIT then it's time for the American people to do a BREXIT.  ""Vote Trump"" https://"
JoeKoffee|JJohnsonLaw|-0.4588|0.303|0.506|0.191|RT @JJohnsonLaw: Trump supporter and Gun in same sentence. Predictably awful results. https://t.co/ebAOW3chHF
JoeKoffee|twitter|-0.4588|0.303|0.506|0.191|RT @JJohnsonLaw: Trump supporter and Gun in same sentence. Predictably awful results. https://t.co/ebAOW3chHF
PEN_dricklamar|TheFunnyVine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
PEN_dricklamar|vine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
JohnReesePOl|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
JohnReesePOl|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
CallmeWunWun|jordan_stratton|0.0|0.0|1.0|0.0|RT @jordan_stratton: Trump's concession speech is going to be 5-7 minutes of him claiming he never ran for president.
JrmezaMeza|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
JrmezaMeza|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
JacksonJoshua73|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
JacksonJoshua73|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
yousuckmuchass|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
Yonce7Twice|hosthetic|-0.2617|0.173|0.656|0.171|"RT @hosthetic: Trump won Kentucky, but is anyone even surprised? all they do there is fuck and marry their cousins anyways."
martinhanratty|jasonvolack|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
martinhanratty|twitter|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
GermyAnd|NorthTampaTrump|0.0|0.0|1.0|0.0|"RT @NorthTampaTrump: #OH #NC #NH will deliver for Trump. #Florida voters, it is all on you now! Get to the polls and stand in line! Close s"
humaneffect|twitter|-0.3595|0.185|0.815|0.0|Hillary NEEDS YOUR VOTE.Trump is getting Indiana.send a message now. no trump! https://t.co/dy4nAUJB06
Brian_Killeen|twitter|-0.2124|0.22|0.551|0.228|Personally...I don't give a damn whether Trump or his evil brood accepts the results. https://t.co/RieUNvb0x9
chrisandm|twitter|0.3521|0.127|0.6|0.274|"Well said, Tommy!  I couldn't agree more!  Forget Clinton &amp; Trump, #ImWithTommy #ElectionDay https://t.co/Oh4165A5fU"
vignettes7642|KGBVeteran|0.0|0.0|1.0|0.0|RT @KGBVeteran: Black man flashes Trump #MAGA hat at camera. This is in Cleveland. #ElectionDay https://t.co/qw0NzwHksv
vignettes7642|twitter|0.0|0.0|1.0|0.0|RT @KGBVeteran: Black man flashes Trump #MAGA hat at camera. This is in Cleveland. #ElectionDay https://t.co/qw0NzwHksv
Lindseycakes|ygselena|-0.5423|0.412|0.588|0.0|RT @ygselena: Fuck Donald Trump  #ElectionNight
mvrleysky|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
mvrleysky|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
IrishSix1|Democrat_4Trump|0.6249|0.0|0.819|0.181|RT @Democrat_4Trump: Poll closing by STATE.Get out and vote if you haven't done so yet. Trump NEEDS EVERY VOTE. We want to win folks. @rea
svogel2|tponews|0.8016|0.0|0.76|0.24|"RT @tponews: Go vote please. If you see an exit pollster, please feel free to tell them you voted for Trump and why! We have to get the wor"
shyannanicole_|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
shyannanicole_|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
Kwadwo_lancelot|br_uk|0.4767|0.0|0.763|0.237|RT @br_uk: Frank Lampard is fascinated by Donald Trump #ElectionDay https://t.co/ob4yyjAfPd
Kwadwo_lancelot|twitter|0.4767|0.0|0.763|0.237|RT @br_uk: Frank Lampard is fascinated by Donald Trump #ElectionDay https://t.co/ob4yyjAfPd
KurtEarl14|CodyCaseNoSpace|0.1872|0.134|0.682|0.184|@CodyCaseNoSpace It sends a message to the Republican Party that Trump isn't acceptable.
ClftnCllns76|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
ClftnCllns76|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
hesthatguy1986|Kimball1Kelly|0.0|0.0|1.0|0.0|"@Kimball1Kelly Kentucky, one of the coal miner states, keeps bouncing back and forth between 68-74 percent Trump."
EllenBWriter|Ronraj777|0.4404|0.0|0.847|0.153|RT @Ronraj777: Exit Poll: Clinton 53% to Trump 42% Clinton +11 Better For Foreign Policy #ImWithHer https://t.co/I3yUwYRgZ2
EllenBWriter|twitter|0.4404|0.0|0.847|0.153|RT @Ronraj777: Exit Poll: Clinton 53% to Trump 42% Clinton +11 Better For Foreign Policy #ImWithHer https://t.co/I3yUwYRgZ2
JohnGilson2|PrisonPlanet|0.0|0.0|1.0|0.0|RT @PrisonPlanet: Votes flipped from Trump to Clinton in Pennsylvania. https://t.co/EBnUDITtOd
JohnGilson2|twitter|0.0|0.0|1.0|0.0|RT @PrisonPlanet: Votes flipped from Trump to Clinton in Pennsylvania. https://t.co/EBnUDITtOd
Lalalavanya8|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
marthawightman|RagnarWeilandt|0.128|0.173|0.628|0.199|RT @RagnarWeilandt: Donald Trump failed to win a single vote from a living US president... #USElection2016
USNCTM|umpire43|0.2023|0.11|0.719|0.171|RT @umpire43: 2 Clinton supporters tried to bully me in line because of my Chemo hookup.Another Clinton supporter came to my aid then he vo
BlayJha|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
BlayJha|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
dmillerwats|juniorsassyrule|0.2732|0.0|0.84|0.16|RT @juniorsassyrule: Trump supporter pepper sprays voter at Florida polling location https://t.co/zhWIGljgtT
dmillerwats|rawstory|0.2732|0.0|0.84|0.16|RT @juniorsassyrule: Trump supporter pepper sprays voter at Florida polling location https://t.co/zhWIGljgtT
randomsweede|Lrihendry|0.3802|0.0|0.874|0.126|RT @Lrihendry: LOOK who just voted for Donald Trump! His biggest fan and unofficial Trump cartoonist #TRUMPTOON  @realDonaldTrump @Kevlar
POOetryman|JonRiley7|0.4404|0.0|0.879|0.121|"RT @JonRiley7: I'm at Trump's star on the Walk of Fame. It's been vandalized so it's covered in wood, surrounded by protesters.#ElectionDa"
CtBrokerRoks|twitter|0.5255|0.0|0.861|0.139|"Notice the MAGA hat? Of course, he inspected the septic system &amp; is a proud small business owner in Ct! Trump is https://t.co/UWEjwbHOsw"
mcuellar|johnolilly|-0.5255|0.328|0.573|0.099|"RT @johnolilly: Damn, okay. Trumps Tears v2.0: Vodka, bitters, Goldschlager (luxury!), muddled with orange peel."
myhorsecowboy|michelleaukamp|0.0|0.0|1.0|0.0|"RT @michelleaukamp: VOTE VOTE #DRAINTHESWAMP Scientific Poll Shows Trump With ""Yuge"" Lead in Swing States https://t.co/i0H9oawmts via @YouT"
myhorsecowboy|linkis|0.0|0.0|1.0|0.0|"RT @michelleaukamp: VOTE VOTE #DRAINTHESWAMP Scientific Poll Shows Trump With ""Yuge"" Lead in Swing States https://t.co/i0H9oawmts via @YouT"
ValisWatson|HispanicsTrump|0.4374|0.0|0.874|0.126|RT @HispanicsTrump: This election is coming down to the wire. Please if you haven't already get out and vote Trump!! #ElectionDay
Riley_green2020|HispanicsTrump|0.6208|0.107|0.659|0.234|RT @HispanicsTrump: My family didn't immigrate to this great county to be taken over by a criminal. Please do your duty and vote for Trump!
ProudfitAsian|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
aura_doree|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
NewCastleNews|cnhipa|-0.4404|0.206|0.794|0.0|RT @cnhipa: Toomey on voting for Trump: 'I struggled with this decision ... it was a tough call.'
mykaela_watkins|Avstvn|-0.1695|0.196|0.804|0.0|"RT @Avstvn: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
jimjrdetore|SpryGuy|-0.296|0.084|0.916|0.0|RT @SpryGuy: The fact that no living US President or First Lady voted for Donald Trump should speak volumes to his unsuitability to the job
elinepomstra|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
N9ZF|TFinn82|0.0258|0.202|0.64|0.158|"@TFinn82 @SMLBound sorry, I've been pretty attentive and I don't recall Trump EVER uttering such lies. Reference?"
amberglows|MOVEFORWARDHUGE|0.0|0.0|1.0|0.0|"RT @MOVEFORWARDHUGE: ""BREAKING VIDEO : Pennsylvania Voting Machines Flipping Votes From Trump to Clinton"" #mustread #feedly https://t.co/3E"
amberglows|t|0.0|0.0|1.0|0.0|"RT @MOVEFORWARDHUGE: ""BREAKING VIDEO : Pennsylvania Voting Machines Flipping Votes From Trump to Clinton"" #mustread #feedly https://t.co/3E"
clperez_eng|AmericasVoice|-0.2023|0.094|0.848|0.058|RT @AmericasVoice: BREAKING: National exit poll number for Latino Voters from @LatinoDecisions: Clinton 79 - Trump 18. New low for GOP. Sam
Melissa_Moyle|DaRealDanBaulch|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
Melissa_Moyle|t|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
DutraGale|KellyannePolls|0.7096|0.0|0.781|0.219|RT @KellyannePolls: Trump Campaign &amp; RNC @Reince hand in glove. This is about GOP elected officials bragging they voted 3rd party or skippe
JDOZIER66|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: If KY holds anywhere near current levels, Trump will outperform polls there by 35 points."
justinamazing1|Bpfillherup|-0.0258|0.167|0.67|0.163|RT @Bpfillherup: Trump winning all the states where the majority of the people fuck their relatives
FlightNemesis|zakwinfield|0.0754|0.183|0.581|0.236|"RT @zakwinfield: So hopefully when I wake, Trump the twat won't be the next American president. Hopefully  #ElectionNight"
SibsMUFC|mcfccentral|-0.5574|0.192|0.76|0.048|@mcfccentral Can anyone seriously see Trump at the UN or going to a poor area thats just been hit by a hurricane? Its laughable
ErnestLamonica|MattGertz|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
ErnestLamonica|twitter|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
CoolsomeXD|TheSuplexCity|0.0|0.0|1.0|0.0|RT @TheSuplexCity: Message to Donald Trump! https://t.co/nSd7K97SGa
CoolsomeXD|twitter|0.0|0.0|1.0|0.0|RT @TheSuplexCity: Message to Donald Trump! https://t.co/nSd7K97SGa
ECVBanana|ABC|0.0|0.0|1.0|0.0|@ABC they kept running out of Orange Clown food color!  ple vote Nov 28th as your overlord commands!https://t.co/7ip7XDo6XX
ECVBanana|businessinsider|0.0|0.0|1.0|0.0|@ABC they kept running out of Orange Clown food color!  ple vote Nov 28th as your overlord commands!https://t.co/7ip7XDo6XX
nochangeplease|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
gtluna1|washingtonpost|0.4588|0.0|0.857|0.143|Does his attys know of Rule 11? The Trump campaign just basically got laughed out of a Nevada courtroom https://t.co/BfQ8Tvx3fO
PhanTheTakeover|EvanEdinger|0.1531|0.242|0.469|0.289|@EvanEdinger if trump wins I'm going to cry
maddieemacc|priscillux|-0.367|0.27|0.522|0.209|RT @priscillux: I don't care if you're a Trump supporter. I respect everyone's opinions. But racism and sexism aren't opinions.
DNJMerica|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
AnnaLinkous|KingKoIbe|-0.2617|0.194|0.674|0.132|RT @KingKoIbe: Voting Trump but sadly America is filled with too many ignorant people who care more about who Beyonc is voting for than th
sharonawesemo|TODAYonline|0.0|0.0|1.0|0.0|RT @TODAYonline: Photo of #DonaldTrump peeking at wife Melania voting goes viral https://t.co/bU2rKcswPR #USElection2016 https://t.co/Kejg1
sharonawesemo|todayonline|0.0|0.0|1.0|0.0|RT @TODAYonline: Photo of #DonaldTrump peeking at wife Melania voting goes viral https://t.co/bU2rKcswPR #USElection2016 https://t.co/Kejg1
Shorty_343|WORLDSTARC0MEDY|0.3612|0.082|0.781|0.138|RT @WORLDSTARC0MEDY: Stop saying if trump wins yall moving out of the country. Stfu yall cant even move outta ya mommas house https://
Shorty_343||0.3612|0.082|0.781|0.138|RT @WORLDSTARC0MEDY: Stop saying if trump wins yall moving out of the country. Stfu yall cant even move outta ya mommas house https://
SickUncleSam|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
RudyStumpo|lisalponder|0.0|0.0|1.0|0.0|RT @lisalponder: #MAGASELFIE We did it!! Women for Trump!!! https://t.co/MMhIXAgEQI
RudyStumpo|twitter|0.0|0.0|1.0|0.0|RT @lisalponder: #MAGASELFIE We did it!! Women for Trump!!! https://t.co/MMhIXAgEQI
carrendaisy|kindcutesteve|-0.296|0.115|0.885|0.0|RT @kindcutesteve: Dana Milbank: Anti-Semitism is no longer an undertone of Trumps campaign. Its the melody#p2 #TNTweeters #USLatinohtt
CORTES4PREZ|LxuiSavage|0.0|0.0|1.0|0.0|RT @LxuiSavage: Trump tryna take all the lil Spanish fum away from a nigga
DeliaEnriquez|_lexabrown|0.5859|0.115|0.573|0.313|"RT @_lexabrown: however, i have no respect for Trump supporters at all. nada. zilch. zero."
4TheTruth2012|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
szabados31|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
realmirokliment|DonaldJTrumpJr|0.8398|0.0|0.69|0.31|"RT @DonaldJTrumpJr: Please watch and share this. Vote now to take back America! ""Freedom is never more than one generation away from exti"
itzgb53J|AdamsFlaFan|-0.7003|0.266|0.734|0.0|RT @AdamsFlaFan: A Nevada judge gave the Trump campaigns voter fraud paranoia the smackdown it deserved https://t.co/z3o2G7aatR via @voxdo
itzgb53J|vox|-0.7003|0.266|0.734|0.0|RT @AdamsFlaFan: A Nevada judge gave the Trump campaigns voter fraud paranoia the smackdown it deserved https://t.co/z3o2G7aatR via @voxdo
truth4ever87|RawStory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
truth4ever87|rawstory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
HollyNiotti|tio2x13|0.0|0.0|1.0|0.0|RT @tio2x13: Florida residents are voting for Trump in RECORD NUMBERS! They are doing everything to get people to the polls! Carry them on
Bcrook21|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Bcrook21|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
bri_bobcat|Flames_Baldwin|0.3612|0.0|0.889|0.111|"RT @Flames_Baldwin: Today I saw a very white woman holding a ""Chinese Americans for Trump"" sign and I dunno man I just feel like the world"
witnessfacts|FrenchForTrump|0.7058|0.0|0.796|0.204|RT @FrenchForTrump: FOR THE FIRST TIME IN MY LIFEAS A FRENCH EXPATRIATEI'M SO PROUD TO CAST MY VOTEFOR DONALD J. TRUMP#ElectionDay#Vo
AscanioMatt|muzikgirl11|0.4084|0.173|0.564|0.263|RT @muzikgirl11: PLEASE everyone who is anxious &amp; fearful. Remember BREXIT. We are having our own BREXIT - AMER-EXIT. Have faith. God will
Amyloukingery|chuckwoolery|0.3182|0.133|0.663|0.204|"RT @chuckwoolery: If #Trump wins, I can't wait to find out who the #Democrats blame."
Captain_Hudson|twitter|0.3612|0.0|0.828|0.172|Trump's cake looks like it just found out it's Trump's cake. #ElectionNight https://t.co/NcOb0RMpo3
GlkEquiped|mitchellvii|0.4404|0.0|0.805|0.195|"RT @mitchellvii: Trump leads IND 72-25.  Good Lord people, something is happening here."
toflyyyyjust|SheHatesJacoby|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
toflyyyyjust|twitter|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
milicopeland|LateNightSeth|0.0|0.0|1.0|0.0|RT @LateNightSeth: From tonights #ACloserLook: How could anyone choose between Trump and Clinton? https://t.co/lUc6pVY3D5
milicopeland|twitter|0.0|0.0|1.0|0.0|RT @LateNightSeth: From tonights #ACloserLook: How could anyone choose between Trump and Clinton? https://t.co/lUc6pVY3D5
FortuneClint|youtube|0.0|0.0|1.0|0.0|Voting machines in Pennsylvania switch Trump votes to Hillary https://t.co/MB4HMHDGbb
amigoalfil|HillaryClinton|0.0772|0.0|0.942|0.058|"RT @HillaryClinton: ""Its not just my name or Donald Trumps name on the ballotits the kind of country we want. Hillary https://t.co/jf"
amigoalfil|t|0.0772|0.0|0.942|0.058|"RT @HillaryClinton: ""Its not just my name or Donald Trumps name on the ballotits the kind of country we want. Hillary https://t.co/jf"
RdzMarisoll|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
FletcherCbpaws|Jpat1952|0.505|0.114|0.676|0.21|RT @Jpat1952: Don't trust ANY polls!!...Go out and vote anyway. We need to give TRUMP a BREXIT win!! https://t.co/BO329Cf2ic
FletcherCbpaws|twitter|0.505|0.114|0.676|0.21|RT @Jpat1952: Don't trust ANY polls!!...Go out and vote anyway. We need to give TRUMP a BREXIT win!! https://t.co/BO329Cf2ic
CharlieEricks10|LarryT1940|0.0|0.0|1.0|0.0|RT @LarryT1940: #Vote4Trump and don't let these #Slime_balls of #Hillary's drive you away from voting. Your vote may push #Trump over the t
KareemLumumba|dailymail|0.0|0.0|1.0|0.0|Trump booed as he votes with Melania and Ivanka in Manhattan https://t.co/sKxCsmFh1G
kanimozhi|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Keylorinho|OdegaardEsque|0.0|0.0|1.0|0.0|RT @OdegaardEsque: Trump masterclass incoming https://t.co/0jxzY3lYSP
Keylorinho|twitter|0.0|0.0|1.0|0.0|RT @OdegaardEsque: Trump masterclass incoming https://t.co/0jxzY3lYSP
Rashaad_DaDon|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Rashaad_DaDon|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
nordicscripts|WordSmithGuy|0.8658|0.0|0.65|0.35|"RT @WordSmithGuy: As a Ted Cruz Constitutional Conservative, I considered who will save the Supreme Court, grow jobs &amp; keep us safe. I vote"
Junkoxxx5|EvanParkerXXX|0.5972|0.0|0.83|0.17|"RT @EvanParkerXXX: Everyone get your asses out &amp; vote!!  (Unless voting for Trump, feel free to stay at home ) https://t.co/HFqzmFbYjm"
Junkoxxx5|twitter|0.5972|0.0|0.83|0.17|"RT @EvanParkerXXX: Everyone get your asses out &amp; vote!!  (Unless voting for Trump, feel free to stay at home ) https://t.co/HFqzmFbYjm"
WhaleLordNorth|ditzkoff|0.0|0.0|1.0|0.0|RT @ditzkoff: Eric Trump gonna Eric Trump https://t.co/JaM3KMhLkL
WhaleLordNorth|twitter|0.0|0.0|1.0|0.0|RT @ditzkoff: Eric Trump gonna Eric Trump https://t.co/JaM3KMhLkL
inukshukuk2|stephenWalt|-0.34|0.098|0.902|0.0|RT @stephenWalt: Imagine being the staffer asked to draft #Trump concession speech (if he intends to make one). How many people can u blame
skepticsmash|DoyleMcManus|0.0|0.0|1.0|0.0|"RT @DoyleMcManus: @AnnCoulter None of Trump's four grandparents were born in the US. Two in Germany, two in UK. A nation of immigrants!"
MarliDivine|RealBenCarson|0.8395|0.0|0.64|0.36|@RealBenCarson I did &amp; I am hoping for Trump/Pence win &amp; U playing a major role in his cabinet! MAGA...Ga in the house!
Mahaksapatalika|Rambobiggs|0.0|0.0|1.0|0.0|"@Rambobiggs Trump, all the way."
diaaanuuuh|SportsTakeJames|-0.1531|0.117|0.789|0.094|RT @SportsTakeJames: Choosing between Hillary &amp; Trump to replace Obama is like when the McDonald's ice cream machine is broken &amp; you gotta
juliann23_|elias_chairez|-0.2348|0.212|0.635|0.153|RT @elias_chairez: People giving Hillary their vote so Trump won't win: https://t.co/0SfLCKj03a
juliann23_|twitter|-0.2348|0.212|0.635|0.153|RT @elias_chairez: People giving Hillary their vote so Trump won't win: https://t.co/0SfLCKj03a
KelliBHorne|Trump2016News|0.0|0.0|1.0|0.0|"RT @Trump2016News: Republicans: I know you're all busy WORKING, but don't put off voting at 5PM! Trump never gave up on you; don't give up"
BeckyMckenzie|PaulbernalUK|-0.5423|0.259|0.741|0.0|RT @PaulbernalUK: I think Trump *can* bring change. All of it bad.
thefridaybarn|JohnKStahlUSA|-0.8519|0.368|0.632|0.0|RT @JohnKStahlUSA: Undocumented relative charged with killing 10-year-old girl. Still think Trump was wrong? #tcot #ccot #gop #maga  https:
ajaimeew|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
ajaimeew|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
heinzman_jo|fightingmajor1|0.2461|0.076|0.81|0.114|RT @fightingmajor1: @mitchellvii If you look at Breibart exit poll headlines it SCREAMS Trump but still who knows for sure. I think it will
vorpalpoet|HeadlineSmasher|-0.5423|0.368|0.632|0.0|RT @HeadlineSmasher: Trump Expected to Destroy Trump
reillyfuller|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
SeanXiao8|0hour|0.0|0.0|1.0|0.0|RT @0hour: Kentucky Trump 69% Lads!
LAMOONLYNN|DiamondandSilk|0.0|0.0|1.0|0.0|"RT @DiamondandSilk: .@realDonaldTrump is Americans only Choice.  Blacks, whites, Hispanics, Asian, Latinos  Vote, Vote, Vote. ......Vote Tr"
AmericanMom2|briojaxen|0.4215|0.1|0.71|0.19|"RT @briojaxen: And if trump looks like winning, they will say its a Russian cyber attack, and you know how that will go. They are already"
Kians_Baddie|ygselena|-0.5423|0.412|0.588|0.0|RT @ygselena: Fuck Donald Trump  #ElectionNight
russmove|mitchellvii|0.5719|0.0|0.85|0.15|"RT @mitchellvii: Romney won Brevard County by 36,000 votes in 2012.  I calculate Trump leads it by 52,000 votes.  +16,000 votes for Trump o"
howell1_howell|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
howell1_howell|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
Kathywa48814788|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
Kathywa48814788|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
__shi_ge__|sharonclott|-0.6249|0.282|0.718|0.0|RT @sharonclott: Protest inside polling station where Trump votes. Two women arrested. #Election2016 #vote https://t.co/YxXKb8NwMD
__shi_ge__|twitter|-0.6249|0.282|0.718|0.0|RT @sharonclott: Protest inside polling station where Trump votes. Two women arrested. #Election2016 #vote https://t.co/YxXKb8NwMD
Azingra76|mitchellvii|0.2177|0.137|0.684|0.179|RT @mitchellvii: So was Trump winning CO and conveniently every voting machine in the state broke?
jayla_laine|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
australian|antfarmer|0.4927|0.0|0.849|0.151|RT @antfarmer: Paul Kelly is very good here on Trump as a vandal and the decline of America ($) https://t.co/ydGRKhuvHc
australian|theaustralian|0.4927|0.0|0.849|0.151|RT @antfarmer: Paul Kelly is very good here on Trump as a vandal and the decline of America ($) https://t.co/ydGRKhuvHc
ElminaNovikova|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ElminaNovikova|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
Hickory_dickery|The_Servant10|-0.3612|0.091|0.909|0.0|RT @The_Servant10: they say the election rigged if trump loses.. same thing my people say when we get pulled over or when we gotta dig anot
fern_friend21|thejournalista|-0.5574|0.247|0.753|0.0|RT @thejournalista: Eric Trump tweets then deletes an illegal ballot selfie. https://t.co/Gjd0aQtlTu
fern_friend21|twitter|-0.5574|0.247|0.753|0.0|RT @thejournalista: Eric Trump tweets then deletes an illegal ballot selfie. https://t.co/Gjd0aQtlTu
SaraKellar|talkwordy|-0.4019|0.13|0.87|0.0|"RT @talkwordy: ""Joe get the Trans Am gassed up we're going to New York to crash Trump's par--"" https://t.co/dUwi0B8QQt"
SaraKellar|twitter|-0.4019|0.13|0.87|0.0|"RT @talkwordy: ""Joe get the Trans Am gassed up we're going to New York to crash Trump's par--"" https://t.co/dUwi0B8QQt"
niki_alisha1|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
niki_alisha1|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
4lovesingaza|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Alex_Derouen|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
RondaBradley00|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
RondaBradley00|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
MataoWilliams|popss0n|0.7003|0.0|0.58|0.42|RT @popss0n: If trump wins I will believe in god again
springspiritual|VladimirPutin24|0.0|0.0|1.0|0.0|RT @VladimirPutin24: Don't Let Donald Trump Put Vladimir Putin in the White House - Heat Street https://t.co/t0hGlFus5a
springspiritual|heatst|0.0|0.0|1.0|0.0|RT @VladimirPutin24: Don't Let Donald Trump Put Vladimir Putin in the White House - Heat Street https://t.co/t0hGlFus5a
KeswickPinhead|SenFallon2016|0.2481|0.089|0.786|0.125|"RT @SenFallon2016: This election is rigged! I intended to vote for #Trump today, when Jesus smacked me upside the head &amp; made my hand vote"
xDrakeFam|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
xDrakeFam|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
LRedderso|halsteadg048|-0.7184|0.222|0.778|0.0|"RT @halsteadg048: Trump Voters, let NOTHING the media says today discourage you.  Make this the LAST time they steal a vote with a lie. htt"
baethompson|twitter|0.4503|0.088|0.716|0.196|"No, they can. Trump tried to sue and so people couldn't but he failed https://t.co/MDlS7tMq7U"
anesiadiego|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
bdarlingwhite|ananavarro|-0.2732|0.087|0.913|0.0|"RT @ananavarro: Hey Nevadans, u know why Trump is suing? To keep Hispanics from polls b/c he knows we're voting against him. Redouble your"
BDChadwick|CKHUK|0.5719|0.0|0.802|0.198|"RT @CKHUK: @BDChadwick if Trump wins and starts WW3, can I be excused from WBAs this year?"
cutestphiI|pastelphilly|-0.5423|0.201|0.712|0.087|RT @pastelphilly: anyways if you support trump at all youre a ignorant shithead in my book dont talk to me &amp; deactivate while youre at it 
charprat44|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
charprat44|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
officiallykumar|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
hibadjedaini|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
BoothRegboo|vandives|0.4753|0.0|0.853|0.147|"RT @vandives: I just voted for our next president, Donald J. Trump  a true American patriot &amp; the ultimate MADMAN!#MAGA3X #MAGASELFIE "
alyssaaafreeman|brooke_hawley5|-0.872|0.319|0.681|0.0|RT @brooke_hawley5: Hmmm  would I rather vote for a woman who helped her rapist husband or a righteous racist in Donald Trump? I'll take D
Voivode_|jackbgoode1|0.0|0.0|1.0|0.0|RT @jackbgoode1: &amp; they vote for this... - VOTE TRUMP @DonaldTrumpVote @USFreedomArmy @Karennola719 @Jnbarke @realDonaldTrump https://t.co/
Voivode_|t|0.0|0.0|1.0|0.0|RT @jackbgoode1: &amp; they vote for this... - VOTE TRUMP @DonaldTrumpVote @USFreedomArmy @Karennola719 @Jnbarke @realDonaldTrump https://t.co/
mltrickey|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
commonsense258|jaynordlinger|0.4404|0.0|0.884|0.116|RT @jaynordlinger: If Bill Clinton talked Donald Trump into running for the GOP nomination -- Clinton truly is the wiliest politician in wo
jnjbowtique|megynkelly|0.0|0.0|1.0|0.0|"RT @megynkelly: 18 electoral votes are up for grabs in #Ohio, and the states own Republican Gov. John Kasich says he did not vote for #Tru"
Worped4|ILoveBernie1|-0.8689|0.329|0.671|0.0|"RT @ILoveBernie1: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, https"
MyNameIsNotMina|Amlx_o|0.4753|0.0|0.808|0.192|"RT @Amlx_o: ""And the next president of the United States is Donald Trump!"" https://t.co/oEIVNItHEE"
MyNameIsNotMina|twitter|0.4753|0.0|0.808|0.192|"RT @Amlx_o: ""And the next president of the United States is Donald Trump!"" https://t.co/oEIVNItHEE"
KatEdmiston|BruceBartlett|0.6311|0.076|0.688|0.235|"RT @BruceBartlett: For the record, I voted enthusiastically for Hillary Clinton today. She may not be perfect, but she's light years better"
ChiefCRX340|BlastingNews|0.0|0.0|1.0|0.0|RT @BlastingNews: #election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR http
ChiefCRX340|us|0.0|0.0|1.0|0.0|RT @BlastingNews: #election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR http
mclvicencio|nytimes|-0.296|0.167|0.833|0.0|"Without Florida, Trump has no path. Polls there close in a minute.  https://t.co/DWteJRFTsB"
Eykis|JRehling|-0.3612|0.116|0.884|0.0|RT @JRehling: Donald Trump started life with a $14 million loan from his father.He thinks the system is rigged against him.#ElectionNight
SteveGoldwing|AMTrump4PRES|0.5255|0.0|0.881|0.119|"RT @AMTrump4PRES: One proud mama hereMy 18 year old son just voted for the first time for the next President of the USA, Donald J. Trump!"
BenShapiro2020|mitchellvii|0.5267|0.0|0.702|0.298|"I heard trump is winning California, can you confirm @mitchellvii ?"
BestWebEnglish|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
70LeRoy|fw|-0.3818|0.205|0.667|0.129|"1 dead, multiple people shot near Azusa polling station; active shooter heavily armed, officials said https://t.co/bTEwV7v6oZ#TRUMP LEGACY"
Magnus_Jamieson|pastachips|0.8658|0.0|0.637|0.363|"@pastachips people with trump avatars and ""deplorable"" in their profiles are liking and sharing it, i am living my best life"
JustMyOwnOpnion|politico|0.0|0.0|1.0|0.0|@politico @PTicks Wasn't the common understanding that not voting works out 2b a vote for Trump?
carsonutt|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Hbb2699|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: 90% of America does not approve of Congress &amp; Washington DC. Trump will DRAIN THE SWAMP! #MAGA
zoombouse|tjhutson|0.4926|0.0|0.715|0.285|RT @tjhutson: @NC5_JasonLamb @mitchellvii @NC5 good news for Trump!
soleileva31|stephstabile8|0.0|0.0|1.0|0.0|RT @stephstabile8: trump &gt; hillary
727times|blackmarvelgirl|-0.3612|0.258|0.569|0.174|"RT @blackmarvelgirl: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost"
The_HighLife23|YFNLUCCl|-0.6408|0.514|0.486|0.0|RT @YFNLUCCl: FUCK DONALD TRUMP.
MUSinfonian|GotHot50|0.6708|0.0|0.807|0.193|@GotHot50 not saying trump is any better but the fact that she hasn't gone to prison for something I know I immediately would be says it all
CmiloseMilose|cnni|0.0|0.0|1.0|0.0|"RT @cnni: What a difference an ""r"" makes: Jake Tapper fact-checks Donald Trump's tweet https://t.co/CROFORgoqE #CNNElection https://t.co/wH"
CmiloseMilose|cnn|0.0|0.0|1.0|0.0|"RT @cnni: What a difference an ""r"" makes: Jake Tapper fact-checks Donald Trump's tweet https://t.co/CROFORgoqE #CNNElection https://t.co/wH"
aNickel4thought|jasonvolack|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
aNickel4thought|twitter|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
franco_dimuro|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
franco_dimuro|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
WaltyAlvarez|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Mariaebrothert2|TawnyaSchultz4|0.508|0.0|0.733|0.267|RT @TawnyaSchultz4: We voted. Yes! Trump WILL be President! https://t.co/YQq7IDukAZ
Mariaebrothert2|twitter|0.508|0.0|0.733|0.267|RT @TawnyaSchultz4: We voted. Yes! Trump WILL be President! https://t.co/YQq7IDukAZ
tlvrp_russia|therussophile|-0.3612|0.143|0.857|0.0|#Moscow #SaintPetersburg Nine Ways the U.S. Voting System Is Rigged But Not Against Donald Trump https://t.co/B9thVprAng
Mrgee_bande|Telegraph|0.0|0.0|1.0|0.0|RT @Telegraph: Florida polls start closing in less than 10 minutes. It's a crucial state to watch on #ElectionNight https://t.co/CJCBsKKKNE
Mrgee_bande|telegraph|0.0|0.0|1.0|0.0|RT @Telegraph: Florida polls start closing in less than 10 minutes. It's a crucial state to watch on #ElectionNight https://t.co/CJCBsKKKNE
Drjoyce54|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
ghostofhypotia|JuddLegum|-0.1027|0.128|0.765|0.107|RT @JuddLegum: Trump black outreach strategy:1. Your lives are miserable2. You have nothing to lose3. Beyonc sucks
alanaarosee|dubstep4dads|0.0|0.0|1.0|0.0|RT @dubstep4dads: trump: what are you drawingmelania: uhh... nothing https://t.co/2EMzgUx8yc
alanaarosee|twitter|0.0|0.0|1.0|0.0|RT @dubstep4dads: trump: what are you drawingmelania: uhh... nothing https://t.co/2EMzgUx8yc
Melly_belly29|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
JimJimbo54|DonaldJTrumpJr|0.0|0.0|1.0|0.0|"@DonaldJTrumpJr add one more for Trump, total from this family 5 votes for Trump HRC 0 all from the state of Pa.Vote Trump"
Filterlbc|AltStreamMedia|0.0258|0.139|0.717|0.143|"RT @AltStreamMedia: Judge to Trump: ""Only you can bring Hillary to justice. Our corrupt judicial system has failed, #LockHerUp"""
INFOS_EN|belfasttelegraph|0.25|0.0|0.824|0.176|US election results: Donald Trump and Hillary Clinton await their verdict of voters - Belfast Telegraph https://t.co/ypMwah7jqC
_Tyreeezy|ciccmaher|0.7738|0.074|0.575|0.351|"RT @ciccmaher: People losing friends over #Clinton vs. #Trump, but guess who's not gonna stop being friends? https://t.co/ctFcxlMEyL"
_Tyreeezy|twitter|0.7738|0.074|0.575|0.351|"RT @ciccmaher: People losing friends over #Clinton vs. #Trump, but guess who's not gonna stop being friends? https://t.co/ctFcxlMEyL"
PrincessJamie47|vnicolesosa123|-0.7378|0.284|0.624|0.092|RT @vnicolesosa123: What gets me mad is seeing latinos with IMMIGRANT PARENTS or FAMILY MEMBERS voting for trump like WTF
RupaStein|Bill_Nye_Tho|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
RupaStein|twitter|0.4404|0.0|0.838|0.162|RT @Bill_Nye_Tho: rt if u think this tiny squid would be a better president than donald trump https://t.co/3zdz5DNTB5
memeswearmatty|letters2donald|0.0|0.0|1.0|0.0|"RT @letters2donald: Children's letters to Donald Trump:  I saw Hilary cheet at hopscotch.Mauvais G., age 8"
CathyMAGA|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
CathyMAGA|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
andywue|laurenasarson|-0.6436|0.239|0.672|0.088|"RT @laurenasarson: The fact that women vote for Trump because ""their husbands talk like that"" is even more disheartening and disgusting. #E"
shonselysees|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
shonselysees|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
ekujpg|jacksfilms|0.0|0.0|1.0|0.0|RT @jacksfilms: You only have a few hours left to write your Trump/Hillary fanfiction
karbripal3|yankeebrit77|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
karbripal3|twitter|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
aeoost|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
aeoost|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
old_put|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
patchrhythm|cyberzlut|0.4019|0.113|0.696|0.192|RT @cyberzlut: WHY IS TRUMP WINNING IM GETTING ANXIETY OVER THIS AND IM NOT EVEN AMERICAN https://t.co/01C70A0bRz
patchrhythm|twitter|0.4019|0.113|0.696|0.192|RT @cyberzlut: WHY IS TRUMP WINNING IM GETTING ANXIETY OVER THIS AND IM NOT EVEN AMERICAN https://t.co/01C70A0bRz
Namndhela|Princessofwifi|-0.3724|0.203|0.797|0.0|RT @Princessofwifi: This is why Donald Trump can't be trusted https://t.co/pmXb95SbLD
Namndhela|twitter|-0.3724|0.203|0.797|0.0|RT @Princessofwifi: This is why Donald Trump can't be trusted https://t.co/pmXb95SbLD
Westxgal|randy_covington|0.4939|0.0|0.802|0.198|RT @randy_covington: @bfraser747 @Westxgal we have to follow through. Save America #MAGA vote #Trump
wtati78|CNN|0.0|0.0|1.0|0.0|"RT @CNN: Ana Navarro: I'm a Republican but voted for Clinton; ""Rather, I cast my vote against Donald Trump"" https://t.co/AN2hI8XFVE via @CN"
wtati78|cnn|0.0|0.0|1.0|0.0|"RT @CNN: Ana Navarro: I'm a Republican but voted for Clinton; ""Rather, I cast my vote against Donald Trump"" https://t.co/AN2hI8XFVE via @CN"
makaylasinspace|keaneyy_|0.5719|0.0|0.829|0.171|RT @keaneyy_: If i wake up and trump's won i'm going back to sleep and not waking up ever again
debbiejoyjoy_|tanamongeau|0.4941|0.0|0.824|0.176|RT @tanamongeau: IF U CAN VOTE fuckin vote !!!! DO U WANT DONALD FUCKING TRUMP AS UR PRESIDENT
wendihoes|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
wendihoes|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
FlySince91_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
FlySince91_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
pattylynn51|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
Bhoysagoodin|RepStones|-0.8908|0.37|0.63|0.0|"RT @RepStones: Trump has more failed businesses and bankruptcies than the rest of Wall Street put together, he's a moron ffs https://t.co/1"
Bhoysagoodin|twitter|-0.8908|0.37|0.63|0.0|"RT @RepStones: Trump has more failed businesses and bankruptcies than the rest of Wall Street put together, he's a moron ffs https://t.co/1"
macariomx|jaynordlinger|0.4404|0.0|0.884|0.116|RT @jaynordlinger: If Bill Clinton talked Donald Trump into running for the GOP nomination -- Clinton truly is the wiliest politician in wo
tom_rowbotham|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
tom_rowbotham|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
doedhavfrue|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
doedhavfrue|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
stacimaione|mitchellvii|0.3182|0.0|0.723|0.277|RT @mitchellvii: Trump leads Kentucky 77-20. :-)
vineandwhimsy|etsy|0.0|0.0|1.0|0.0|Check out this item in my Etsy shop https://t.co/flMvLy2o6G #trump #TrumpPence16 #Election2016 #MAGA #etsy #deplorable
kenD0LLnbarbie|totalfratmove|0.3612|0.0|0.828|0.172|RT @totalfratmove: This Cake Shaped Like Trumps Head Is Nightmare Fuel: https://t.co/CN3yDoVFBK https://t.co/T68VcxfTfL
kenD0LLnbarbie|totalfratmove|0.3612|0.0|0.828|0.172|RT @totalfratmove: This Cake Shaped Like Trumps Head Is Nightmare Fuel: https://t.co/CN3yDoVFBK https://t.co/T68VcxfTfL
jamesbott007|rnlisa64|0.0|0.0|1.0|0.0|RT @rnlisa64: Voted Trump!!! #MAGA https://t.co/FTWASnfuRJ
jamesbott007|twitter|0.0|0.0|1.0|0.0|RT @rnlisa64: Voted Trump!!! #MAGA https://t.co/FTWASnfuRJ
lph20|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
SouthernFlag88|PoliticsWolf|0.0|0.0|1.0|0.0|"RT @PoliticsWolf: Elliott County KY has literally always voted Democratic, even back to the 1820s &amp; before it was formed in the 1860s. Trum"
adafocobo|syoka68|-0.2462|0.099|0.901|0.0|RT @syoka68: Not hard to believe they are rigging exit polls! Turn off the tv GO VOTE TRUMP! https://t.co/HLNXmSp0IQ
adafocobo|twitter|-0.2462|0.099|0.901|0.0|RT @syoka68: Not hard to believe they are rigging exit polls! Turn off the tv GO VOTE TRUMP! https://t.co/HLNXmSp0IQ
StephsterStarrO|NestorMendoza66|0.5696|0.0|0.822|0.178|RT @NestorMendoza66: I'm proud! That my first vote as an American Citizen was for Trump! #MAGASELFIE #MAGA3X https://t.co/kzX5QWCl6M
StephsterStarrO|twitter|0.5696|0.0|0.822|0.178|RT @NestorMendoza66: I'm proud! That my first vote as an American Citizen was for Trump! #MAGASELFIE #MAGA3X https://t.co/kzX5QWCl6M
Bella2169Molina|mitchellvii|0.34|0.0|0.893|0.107|"RT @mitchellvii: I expect Trump to win KY and IN, but not by 50 points.  We'll see if anything near that holds."
magicimpact|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
magicimpact|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
kuhar_l|NewtTrump|0.8866|0.0|0.668|0.332|"RT @NewtTrump: AWESOME: Tom Brady endorses Trump and the crowd in New Hampshire goes WILD! To make it better, Pats Coach Bill Belichick als"
angxlxsxphxa|VictoriaAveyard|0.7269|0.136|0.568|0.297|"RT @VictoriaAveyard: ""It would be sweet sweet justice if it was the Latino vote that stopped Trump."" - Ana Navarro continuing to spit fire."
anahi__16|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
anahi__16|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
Politicalife|francishumes|0.0|0.0|1.0|0.0|RT @francishumes: Spent my lunch hour dropping off our ballots and stumping for Trump! The Cappello's have officially voted for @realDonald
not_prescott|RowdyAmericans|0.0|0.0|1.0|0.0|RT @RowdyAmericans: Now that all the Republicans are off work it's time to Trump the polls
jewelbird918|TheTylt|0.3182|0.122|0.667|0.212|RT @TheTylt: RT if you agree Ivanka Trump ruined her own brand by supporting her misogynist father #IvankaIsToast #BoycottIvanka https://t.
jewelbird918||0.3182|0.122|0.667|0.212|RT @TheTylt: RT if you agree Ivanka Trump ruined her own brand by supporting her misogynist father #IvankaIsToast #BoycottIvanka https://t.
betteranfiction|shootist2015|0.0|0.0|1.0|0.0|RT @shootist2015: #Florida we can't do this without you.  Get out there and cast that vote for #Trump for change and to #MAGA and #drainthe
CKlein5852|AdamsFlaFan|0.0|0.0|1.0|0.0|RT @AdamsFlaFan: Hillary Clinton Is Trouncing Trump With Her Ground Game According To Exit Poll via @politicususa https://t.co/Fa8OqrLYog
CKlein5852|politicususa|0.0|0.0|1.0|0.0|RT @AdamsFlaFan: Hillary Clinton Is Trouncing Trump With Her Ground Game According To Exit Poll via @politicususa https://t.co/Fa8OqrLYog
Waja1130|kmbiamnozie|0.0|0.0|1.0|0.0|"RT @kmbiamnozie: An estimated 150,000 Haitian-American voters live in Florida, the state where 537 votes decided the 2000 election, Trump"
kateloving|ErikH526|0.6467|0.0|0.799|0.201|"RT @ErikH526: Watch the latest @HAGOODMANAUTHOR segment!!WIKILEAKS 1-35 BREAKING NEWS: Donald Trump Wins Florida, OH, NC Despite Clinton M"
Clarembaldo|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
Carinamarie123|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
PatriotesLibres|DonaldJTrumpJr|0.8279|0.079|0.638|0.283|RT @DonaldJTrumpJr: Freedom is never more than one generation away from extinction. My father will fight for YOU! He will WIN FOR YOU! #Tru
Utdmariam|hucks6dh6|0.807|0.0|0.735|0.265|"RT @hucks6dh6: Good people of America, please don't vote in Trump, how could this end be in control of the most powerful country in the Wo"
sophia_bonoma|BruhhhComedy|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
sophia_bonoma|twitter|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
africanvodka|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
ChuckCollier76|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @MaddieAndMichi @enjoynChi @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE
leidasavina87|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
leidasavina87|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
Suave_young50|twitter|0.3612|0.0|0.615|0.385|You look like trump https://t.co/UYplEJoKGK
kphbritt|buzzfeed18|0.0|0.0|1.0|0.0|RT @buzzfeed18: Ivanka Trumps poise and polish artfully mask just how closely her ideologies align with her fathers. https://t.co/2cTbpFR
kphbritt|t|0.0|0.0|1.0|0.0|RT @buzzfeed18: Ivanka Trumps poise and polish artfully mask just how closely her ideologies align with her fathers. https://t.co/2cTbpFR
nancymarie4159|BinsackSb|-0.6981|0.243|0.757|0.0|RT @BinsackSb: AMERICA STAND UP NOW!! #DonaldTrump announces lawsuit against Nevada for poll workers wearing defeat Trump T Shirts! Make th
volpappaw|mike_pence|0.4926|0.0|0.849|0.151|RT @mike_pence: Trump Force 2 has landed in NYC! Thanks to everyone who has joined us on this journey. https://t.co/PRaQcEME2G
volpappaw|twitter|0.4926|0.0|0.849|0.151|RT @mike_pence: Trump Force 2 has landed in NYC! Thanks to everyone who has joined us on this journey. https://t.co/PRaQcEME2G
insomniaclucas|EvanEdinger|0.0258|0.281|0.36|0.36|@EvanEdinger trump won kentucky and i want to die
linnyitssn|TeaPartyCat|-0.547|0.22|0.714|0.066|"RT @TeaPartyCat: It's not fair to call all Trump's supporters racist and sexist. Some are racist, some are sexist, but not all of them are"
tnelson027|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
tnelson027|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
michellet0624|Aaronjackson81|0.3612|0.0|0.902|0.098|RT @Aaronjackson81: I like how the news is saying nothing about the voting machines are not allowing  trump voters to vote for trump in swi
dominicxsmith|freeskimask45|0.1258|0.17|0.596|0.234|"@freeskimask45 I would like an answer to my question, so please, tell me how Donald Trump is a racist."
JanelleMonae|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
JanelleMonae|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
ejoy2270|XCrvene|0.4404|0.0|0.888|0.112|"RT @XCrvene: Reports are turn out in the Florida panhandle is under performing. All GOP &amp; Trump supporters in the panhandle, vote Trump now"
KarolineMarquis|BruhhhComedy|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
KarolineMarquis|twitter|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
SexMyTatts|SheHatesJacoby|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
SexMyTatts|twitter|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
chrisg_769|SQUlDZ|0.6841|0.0|0.832|0.168|"RT @SQUlDZ: Mexicans and Black People teaming up against Donald Trump BOY LIFE BEAUTIFUL RN MY NIGGA, bout time tacos and fried chicken uni"
noahtash101|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
noahtash101|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
CS_Perez10|monotonecunt|-0.5423|0.137|0.863|0.0|"RT @monotonecunt: Props to Trump for revealing all of the closet racists, homophobes, sexist &amp; misogynists.. and for showing me who not to"
kaayyrista|Andrea_o0|-0.0516|0.118|0.882|0.0|@Andrea_o0 dude all the old people are for trump i swear
RJC624|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
RJC624|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
pau2la057328721|manusartorius02|-0.5106|0.524|0.476|0.0|RT @manusartorius02: Trump dumb
l_cisneros9|utsafree|0.0|0.0|1.0|0.0|"RT @utsafree: ""I'm voting for Donald Trump!""""why?""""because he's pro-life!""""and?""""that's it!""""wait what?"""
RonaldMRivera|Boogie2988|-0.4019|0.172|0.828|0.0|RT @Boogie2988: Donald trump and Hillary clinton are both in a plane crash.  Who survives?....america.
PurpleRainQuin|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
WinOrGoHome|Only__Trump|0.3802|0.0|0.755|0.245|RT @Only__Trump: @PhillyGOP Vote Trump again &amp; again please!
DTharp1988|FoxNews|0.0|0.0|1.0|0.0|@FoxNews Some will vote for Hillary. Some will vote for Trump. Some will vote AGAINST Hillary or against Trump. I voted for my son's future.
Willsdarlin|BellaSiena|0.6981|0.0|0.781|0.219|RT @BellaSiena: Super long lines in Imperial Pennsylvania. Everyone I talked to was voting for Donald Trump!!! #myvote2016 #ElectionDay2016
realSpottswoode|GartrellLinda|0.2714|0.0|0.905|0.095|RT @GartrellLinda: Important! RTGET OUT THERE &amp; VOTE TRUMPSTERSVERY TIGHT in Florida panhandle. Call everyone you know to get those Trump
Michaelcraddo16|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Michelle3wits|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
Michelle3wits|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
humdinger41|KellyannePolls|0.7096|0.0|0.781|0.219|RT @KellyannePolls: Trump Campaign &amp; RNC @Reince hand in glove. This is about GOP elected officials bragging they voted 3rd party or skippe
WonderLavi|NickKristof|0.0|0.0|1.0|0.0|"RT @NickKristof: But, Anne, then Trump wouldn't vote, because 3 of his 4 grandparents were born abroad, along with his mom. The immigrants"
peachgrI|pupbasket|0.5719|0.0|0.821|0.179|RT @pupbasket: If Trump   Wins The Election I Am Moving   Out Of The Country  Goodbye   America   Hello   EXO Planet 
ocularnervosa|twitter|0.0|0.0|1.0|0.0|In case you donated to Trump's campaign &amp; wondered where the money went. https://t.co/xhFvkOqDNr
an_gonzalez22|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
AnonymousMsBig|SMShow|-0.3818|0.316|0.517|0.167|#Trump supporters blocking polls &amp; intimidating in #Florida@SMShow @frangeladuo @hippiemama2002 @Lawrence https://t.co/sL52VXopWc
AnonymousMsBig|twitter|-0.3818|0.316|0.517|0.167|#Trump supporters blocking polls &amp; intimidating in #Florida@SMShow @frangeladuo @hippiemama2002 @Lawrence https://t.co/sL52VXopWc
mikenziFitz|geena1017|0.3178|0.129|0.697|0.174|@geena1017 well it's a good thing i'm not trying to convince you to vote for trump. i'm just saying he's not responsible for deaths or
fredakalina|thegatewaypundit|-0.4588|0.231|0.769|0.0|Nevada Poll Workers Break Law: Caught Wearing 'Defeat Trump' T-Shirts https://t.co/934mTzlCvd
WillRowland7|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
lemonyspiffit|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
kimmurphy|latimes|0.0|0.0|1.0|0.0|Exit polls: white college-educated voters trending more Democrat than 2012. Non-college educated whites? Trump town. https://t.co/u0nbNhr8ee
HamannRandal|mitchellvii|0.4404|0.0|0.838|0.162|"RT @mitchellvii: If Trump ends up dramatically outperfroming his RCP averages in early states, good sign."
MEAspencer|ananavarro|-0.2732|0.087|0.913|0.0|"RT @ananavarro: Hey Nevadans, u know why Trump is suing? To keep Hispanics from polls b/c he knows we're voting against him. Redouble your"
Zhepon|TeamTrump|0.5781|0.0|0.8|0.2|@TeamTrump @AC360 @ananavarro nice way to talk!lady you mean #Trump woman voters didn't go to college!?Insulating?
francesca281|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
HotlineJosh|NKingofDC|-0.128|0.061|0.939|0.0|"RT @NKingofDC: So far, digging through the exits, and with the first polls about to close, there aren't a lot of signs of a looming Trump u"
kwhunter|twitter|0.3214|0.0|0.795|0.205|"I didn't vote for Trump either, so I don't blame them. https://t.co/4r7qAe5MMj"
melofidias|JaredWyand|0.5859|0.128|0.667|0.206|RT @JaredWyand: It's simple...Trump needs NHIf he loses FL he needs PA &amp; MIIf he wins FL loses NC he needs MI or PAIf he wins FL he
deluxemami|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
deluxemami|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
2babyblueeyes|Madmaven|-0.296|0.216|0.784|0.0|"RT @Madmaven: Say No to Satan, vote TRUMP https://t.co/Y9gulyxgDY"
2babyblueeyes|twitter|-0.296|0.216|0.784|0.0|"RT @Madmaven: Say No to Satan, vote TRUMP https://t.co/Y9gulyxgDY"
DonaldDrumpfWTF|FaithRubPol|-0.296|0.101|0.847|0.052|RT @FaithRubPol: After being criticized for being just a casino promoter that will tell you what you want to hear Trump releases plan https
Artco77|OwensboroMI|0.0|0.0|1.0|0.0|RT @OwensboroMI: With 5 percent of the Kentucky votes in Trump leads by 41 percent.
50shadesofjenny|RAY_2_YAH|0.1999|0.111|0.736|0.153|RT @RAY_2_YAH: The way Donald trump in the lead it don't look like we got hope 
shazzjonz|kurteichenwald|-0.4033|0.244|0.609|0.147|"RT @kurteichenwald: I just realized: With Nevada, Trump is essentially arguing that allowing people to vote is voter fraud. Quite amazing w"
irishowens96|WeLoveRobDyrdek|0.4404|0.0|0.791|0.209|RT @WeLoveRobDyrdek: Jon Stewart and Donald Trump beef is funny af https://t.co/j1HsilMOlH
irishowens96|twitter|0.4404|0.0|0.791|0.209|RT @WeLoveRobDyrdek: Jon Stewart and Donald Trump beef is funny af https://t.co/j1HsilMOlH
sorryimspencerr|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Suweetpea|FredZeppelin12|0.25|0.0|0.895|0.105|RT @FredZeppelin12: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERS. Advantage #Trump. Evening voters are evening voters because t
xoC_Lianne|TomiLahren|0.4717|0.0|0.861|0.139|RT @TomiLahren: If you're not voting for Trump don't you dare bitch when we get Hillary. Real talk. #MAGA #ElectionDay
Women4T|writerkev|0.2732|0.0|0.87|0.13|RT @writerkev: Trump supporter working corner of 120th Avenue and Washington Street. #9NEWS #verifyvotes https://t.co/BVVPseQ1qp
Women4T|twitter|0.2732|0.0|0.87|0.13|RT @writerkev: Trump supporter working corner of 120th Avenue and Washington Street. #9NEWS #verifyvotes https://t.co/BVVPseQ1qp
scooterdawg|krystalball|-0.5267|0.167|0.833|0.0|RT @krystalball: Homes without Trump signs reportedly getting these threatening KKK fliers in rural Kentucky. In 2016. https://t.co/LAGVNbm
scooterdawg|t|-0.5267|0.167|0.833|0.0|RT @krystalball: Homes without Trump signs reportedly getting these threatening KKK fliers in rural Kentucky. In 2016. https://t.co/LAGVNbm
ellawest_|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
CamilleKoch|richthekid|-0.5848|0.256|0.744|0.0|RT @richthekid: If you voting for trump fuck you unfollow me now!
nickgourevitch|NKingofDC|-0.128|0.061|0.939|0.0|"RT @NKingofDC: So far, digging through the exits, and with the first polls about to close, there aren't a lot of signs of a looming Trump u"
DennisL656|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
animalvore|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
Rollo87|Cain_Unable|0.0|0.0|1.0|0.0|"RT @Cain_Unable: I just tried to Vote Trump &amp; the staff wouldn't let me just because I'm ""in Kent"" &amp; ""this is a Tesco self service checkout"
DejaFields127|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
DejaFields127|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
Gyggy|MattGertz|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
Gyggy|twitter|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
KitsuneMonster|Simpsons_tweets|-0.5423|0.163|0.837|0.0|"RT @Simpsons_tweets: ""We've inherited quite a budget crunch from President Trump. How bad is it, Secretary Van Houten?""""We're broke."" #Ele"
PBurgrealtor|kayleighmcenany|0.7177|0.0|0.769|0.231|"RT @kayleighmcenany: Trump has a .2% lead in Florida according to Real Clear Politics. My fellow Floridians, get out, vote, &amp; take friends!"
MelissaBarton|bobcesca_go|-0.2263|0.094|0.851|0.055|RT @bobcesca_go: Here's what I want to see: Khizr Khan interrupting Trump's concession to finally give him his copy of the Constitution. #E
cutebutthood|brujaaverde|-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
cutebutthood||-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
kyotojoe1|abcnews|0.2023|0.0|0.833|0.167|@abcnews @JohnBarronUSA over playing the devil's advocate for Trump? #auspol
Vxwxg33ZsGp6i6I|TommTommmm|-0.5994|0.257|0.632|0.112|@TommTommmm No I am not referring 2 Trump.Clinton just because its a woman one need's to stand on principle non acceptance of rape.
EyasHolden|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
TechL0G|yahoo|0.0|0.0|1.0|0.0|"Trump, the Autocrat's Preferred Choice (Yahoo Security) https://t.co/oKWiSXp8S5"
cryingdun|EvanEdinger|0.7351|0.0|0.53|0.47|@EvanEdinger trump is winning popular vote by quite a bit
dmrider|VassyKapelos|0.0|0.0|1.0|0.0|RT @VassyKapelos: Pro-Trump group in midtown Manhattan https://t.co/dXpgwRJ1BG
dmrider|twitter|0.0|0.0|1.0|0.0|RT @VassyKapelos: Pro-Trump group in midtown Manhattan https://t.co/dXpgwRJ1BG
DjKiddeNJ|ViraI|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
DjKiddeNJ|twitter|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
salngvyen|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
salngvyen|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
leamjavier_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Andrew_Tuft|TBNSport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
Andrew_Tuft|tbnsport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
tiagommmanso|FansOfSport|0.0|0.0|1.0|0.0|RT @FansOfSport: McGregor vs. Trump. #Election2016 https://t.co/2i56Dr4Hlg
tiagommmanso|twitter|0.0|0.0|1.0|0.0|RT @FansOfSport: McGregor vs. Trump. #Election2016 https://t.co/2i56Dr4Hlg
___sunshineee|iEnjoyThoak_DMG|-0.6088|0.312|0.561|0.126|RT @iEnjoyThoak_DMG: I'm bouta get Dronk Dronk hopefully trump don't win and blow my shit
idklife348|ridevocals|-0.4588|0.146|0.778|0.075|"RT @ridevocals: WHY ARE PEOPLE VOTING TRUMP BECAUSE ""HILLARY IS A CRIMINAL"" WHEN THE FBI ALREADY CLEARED HER AND TRUMP IS GOING TO COURT FO"
JDisjuicy|RonnieFieg|0.5719|0.0|0.764|0.236|"RT @RonnieFieg: If Trump wins, going to relocate the team to Kith Canada."
Herfarm|umpire43|0.2023|0.11|0.719|0.171|RT @umpire43: 2 Clinton supporters tried to bully me in line because of my Chemo hookup.Another Clinton supporter came to my aid then he vo
KimberlyFergus|jackbgoode1|0.0|0.0|1.0|0.0|RT @jackbgoode1: Bama's a chimp or is it chump - VOTE TRUMP @DonaldTrumpVote @USFreedomArmy @Karennola719 @Jnbarke @realDonaldTrump https:/
KimberlyFergus||0.0|0.0|1.0|0.0|RT @jackbgoode1: Bama's a chimp or is it chump - VOTE TRUMP @DonaldTrumpVote @USFreedomArmy @Karennola719 @Jnbarke @realDonaldTrump https:/
luisvguevara|Fusion|-0.128|0.113|0.795|0.092|"RT @Fusion: ""Since he's gonna lose, I'm going to go dancing.""Latinas share #ElectionNight predictions at the Nevada store Trump tried &amp; f"
leontiiisaev2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
leontiiisaev2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
HvaMedical|NorthTampaTrump|0.0|0.0|1.0|0.0|"RT @NorthTampaTrump: Folks who just put in a 10 hour shift, u have 5 minutes 2 get in line and vote #trump they can't turn u away if u get"
RAINDROPDOLANS|harrysdolan|0.0|0.0|1.0|0.0|RT @harrysdolan: #ElectionNight what if trump gets elected and the first couple of weeks he's president he gets assassinated LMFAOO
allnighttom|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
HateThisAt|aprendiztg|-0.2032|0.25|0.556|0.194|RT @aprendiztg: donald trump? more like donald DUMP am i right
TeamGOATface|SlackGod|0.0|0.0|1.0|0.0|@SlackGod only reason i voted trump tbh
SamMcCadams|deray|-0.5106|0.125|0.875|0.0|"RT @deray: The @NYTimes has printed a list of all of the people, places, &amp; things that Trump has insulted on Twitter during the campaign. h"
ScottJF666|ScottJF666|0.0|0.0|1.0|0.0|"RT @ScottJF666: Why Why Do they keep saying ""the Non-college white people are voting Republican Trump"" ...?"
raiderfan2466|AlysiaStern|-0.5553|0.146|0.854|0.0|"RT @AlysiaStern: @ananavarro My Hispanic family voted for TRUMP! You don't represent us, in fact you don't REPRESENT. Great work keeping yo"
IsYouMadOrAngry|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
IsYouMadOrAngry|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
Eag1e0ne|MarkDice|-0.4738|0.118|0.882|0.0|RT @MarkDice: Do Hillary voters have to fill out their ballots in blood?  Vote for Trump and let's send that witch into retirement!! #Elect
MOSESMAKASl|georgejxnes|0.0|0.0|1.0|0.0|"@georgejxnes rising sea level London city will be underwater in 100 years, did it in geog, trump doesn't believe in it tho"
andregreen0|CNN|0.6369|0.0|0.833|0.167|"RT @CNN: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/QurbNzL1BK"
andregreen0|cnn|0.6369|0.0|0.833|0.167|"RT @CNN: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/QurbNzL1BK"
njoanyork|PamelaGeller|0.0|0.0|1.0|0.0|"RT @PamelaGeller: Wikileaks: 8,263 NEW emails shows Democrats helped CNN anchors for Trump interviews https://t.co/ppKJgwvtbd"
njoanyork|pamelageller|0.0|0.0|1.0|0.0|"RT @PamelaGeller: Wikileaks: 8,263 NEW emails shows Democrats helped CNN anchors for Trump interviews https://t.co/ppKJgwvtbd"
insomniacsprm|TheDeploring|0.4215|0.0|0.714|0.286|"@TheDeploring true ""*trump is literally the next Hitler"
NotcoolOToole|TheTrumpPuppet|0.0|0.0|1.0|0.0|"RT @TheTrumpPuppet: ""Hello Hillary. How are you doing?"" #Trump #TheTrumpPuppet #Election #ElectionDay https://t.co/iPeB6nFXbl"
NotcoolOToole|vine|0.0|0.0|1.0|0.0|"RT @TheTrumpPuppet: ""Hello Hillary. How are you doing?"" #Trump #TheTrumpPuppet #Election #ElectionDay https://t.co/iPeB6nFXbl"
Richard_RSC|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
Richard_RSC|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
SculptNewYork|KellyannePolls|0.7096|0.0|0.781|0.219|RT @KellyannePolls: Trump Campaign &amp; RNC @Reince hand in glove. This is about GOP elected officials bragging they voted 3rd party or skippe
clanton_jim|twitter|0.0|0.0|1.0|0.0|#Mexicans4 Trump #ElectionNight https://t.co/sTwkHYCUAd
HIGHLYBISEXUAL|THOTJAI|0.5719|0.0|0.821|0.179|RT @THOTJAI: if donald trump wins the election I will paypal 100 dollars to everyone that retweets this #ElectionDay
veeemariee_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
veeemariee_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
scottthong|mitchellvii|0.7227|0.0|0.82|0.18|"RT @mitchellvii: You are leaving out Trump's 5000 vote lead with Indies, so 22,000, but Obama won it by 36,000.  HRC 14,000 behind Obama. h"
Ih8heels|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
pacsgirl36|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
Leandra_C_Lee|lntroset|0.8969|0.0|0.67|0.33|RT @lntroset: Today is Election Day so I thought I would share the loving someone lyrics with you guys bc this world needs more love and le
ThePissBaby|twitter|0.0|0.0|1.0|0.0|Coming to the realization that trump is way ahead in a few states https://t.co/NhRrCF92Ef
Refinery29|refinery29|0.4588|0.0|0.75|0.25|How your favorite celebs are voting during #ElectionDay: https://t.co/OWRZ0dyO0m https://t.co/OyC6vTclZ9
confusednyy|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
confusednyy|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
jihhoons|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
williamcreedcox|vitweet|0.0|0.0|1.0|0.0|CO Voters We Need Your VotesPlease don't do anything after work except VOTE TRUMP! Get to your  #DrainTheSwamp https://t.co/WK9wrWo9gc
NinaaaPadilla|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
NinaaaPadilla|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
HansonbooRiah|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
KayleeGould|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
KayleeGould|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
AuburnFox11|Bencjacobs|0.0|0.0|1.0|0.0|RT @Bencjacobs: Cash bar at trump election night event
sirdrano|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: 90% of America does not approve of Congress &amp; Washington DC. Trump will DRAIN THE SWAMP! #MAGA
balthsbart|twitter|-0.4588|0.234|0.656|0.111|"My Pap was a lifelong #Republican. He would be disgusted beyond words by trumpHe fought nazis, nazis now support t https://t.co/ciwBliRrVP"
2megzzzzz|nrherzog|-0.0258|0.149|0.664|0.187|RT @nrherzog: everyone out here makin' kanye 2020 jokes like shit that's literally how donald trump decided to run
heyit_thatboy|shep689|0.0|0.0|1.0|0.0|RT @shep689: donald trumpdonal trum dona tru don trdont don'tjust don't
kleegrubaugh|KatyTurNBC|-0.4767|0.279|0.721|0.0|@KatyTurNBC @lifebythecreek @chucktodd I am disappointed Trump did not self-fund.
idea15webdesign|seansrussiablog|-0.4939|0.167|0.833|0.0|RT @seansrussiablog: From @GazetaRu live feed. Trump's voting violation hotline. Dial 1 if you're calling from Russia. https://t.co/P12NTVC
idea15webdesign|t|-0.4939|0.167|0.833|0.0|RT @seansrussiablog: From @GazetaRu live feed. Trump's voting violation hotline. Dial 1 if you're calling from Russia. https://t.co/P12NTVC
AFZ33N|Democrat_4Trump|0.6249|0.0|0.819|0.181|RT @Democrat_4Trump: Poll closing by STATE.Get out and vote if you haven't done so yet. Trump NEEDS EVERY VOTE. We want to win folks. @rea
that1BlackGirl|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
that1BlackGirl|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
jrwsjs|recordonline|0.4404|0.0|0.847|0.153|RT @recordonline: Here's what Trump and Clinton supporters are saying about this historic Election Night https://t.co/lgWpBu129k https://t.
jrwsjs|recordonline|0.4404|0.0|0.847|0.153|RT @recordonline: Here's what Trump and Clinton supporters are saying about this historic Election Night https://t.co/lgWpBu129k https://t.
danmthatlady|alkhatib_assil|0.2023|0.0|0.927|0.073|"RT @alkhatib_assil: Muslims or Arabs voting for either Clinton or trump are playing them self, one wants you deported and one wants you kil"
fluffynutters|TrumpDynastyUSA|0.6514|0.0|0.776|0.224|RT @TrumpDynastyUSA: .@realDonaldTrump#TRUMP PULLS the PLUG on DCSay BUH BYE to your FREE RIDE!#DrainTheSwamp #DeplorablePlugPullers #T
joe_bayside|mitchellvii|-0.6186|0.336|0.664|0.0|@mitchellvii BILL FOX IS ALL BUT SAYING TRUMP LOST.
mulasniper|ItsSimplyBeka_3|0.0|0.0|1.0|0.0|@ItsSimplyBeka_3 we just need trump to come through
couchycraig|MagicRoyalty|0.3252|0.059|0.818|0.123|"RT @MagicRoyalty: Hillary doesn't want to #MAGA -- This makes Pepe sad.Please don't make Pepe sad, vote Trump.#ElectionDay https://t.c"
couchycraig||0.3252|0.059|0.818|0.123|"RT @MagicRoyalty: Hillary doesn't want to #MAGA -- This makes Pepe sad.Please don't make Pepe sad, vote Trump.#ElectionDay https://t.c"
BureenuhDuhh|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
BureenuhDuhh|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
legit_leah|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
RobbieBurroughs|kirstiealley|-0.5423|0.2|0.8|0.0|RT @kirstiealley: CELEBS (including myself) R not financially middle or lower M class. U live the bleed. UR $ despair is real. U are being
smelllikesugar|NateMonroeTU|-0.4767|0.134|0.866|0.0|RT @NateMonroeTU: You contrarians are focusing on the wrong thing. It's not whether Trump outperforms '12. It's whether that's enough. May
GoldFramed_|SkyeAsiyanbi|0.3612|0.0|0.872|0.128|RT @SkyeAsiyanbi: If you're voting for Trump today I would like nothing more than for you to unfollow me
BillKS1|DonaldJTrumpJr|0.5696|0.0|0.872|0.128|"RT @DonaldJTrumpJr: If you have friends in MI, OH, FL, PA -- CALL THEM and tell them to VOTE TRUMP! You can make a difference! #MAGA #Tru"
klarolinebonkai|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
klarolinebonkai|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
trumpquility1|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
phil94SR|jeremyscahill|0.6249|0.0|0.661|0.339|RT @jeremyscahill: Trump's final tv ad is a masterpiece: https://t.co/DQK1ZIajP1
phil94SR|twitter|0.6249|0.0|0.661|0.339|RT @jeremyscahill: Trump's final tv ad is a masterpiece: https://t.co/DQK1ZIajP1
GlobeRetroh|RedBeardMLG|0.7579|0.128|0.468|0.404|@RedBeardMLG HRC supporters will keep attacking trump supporters if she wins *cough* rigs it *coughs*
AlicePolidoro|surfermom77|0.0|0.0|1.0|0.0|"RT @surfermom77: Twitter &amp; FB R begin inundated wt reports of Elec.fraud, voting irregularities &amp; discrimination against Trump Votershttps"
FTD_Guido24|sarahmlauren|0.0|0.0|1.0|0.0|"RT @sarahmlauren: President #Trump, it's on the tip of my tongue baby!!! Get out and vote!!! #TrumpPence16 #Trump2016 #TrumpTrain #MakeAmer"
DiRealLauren|megynkelly|0.0|0.0|1.0|0.0|"RT @megynkelly: 18 electoral votes are up for grabs in #Ohio, and the states own Republican Gov. John Kasich says he did not vote for #Tru"
WandaAlbright1|TallahForTrump|0.765|0.0|0.761|0.239|"RT @TallahForTrump: To me, Donald Trump is like a mix between Martin Luther King Jr, Abraham Lincoln, and Cyrus the Great who rebuilt the T"
DeathToAllThots|WhoadieBrees|-0.4003|0.152|0.848|0.0|RT @WhoadieBrees: Niggas with white gfs RT @lovemeGabbi: Who is this 8% voting for trump?! https://t.co/qsNsQ3stvV
DeathToAllThots|twitter|-0.4003|0.152|0.848|0.0|RT @WhoadieBrees: Niggas with white gfs RT @lovemeGabbi: Who is this 8% voting for trump?! https://t.co/qsNsQ3stvV
SlavichMadi|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
SlavichMadi|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
rosetaddie|LaziestCanine|-0.1695|0.196|0.804|0.0|"RT @LaziestCanine: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
shadymendes|s_mxndes|0.8271|0.091|0.514|0.395|RT @s_mxndes: if trump wins can we just hope that kayne west interrupts his winning speech #ElectionNight
sylrei63|mitchellvii|-0.8537|0.377|0.555|0.068|@mitchellvii yes but what counties worried about Date and Broward also low turnout in PanHandleis bad news for Trump
phiI94|jeremyscahill|0.6249|0.0|0.661|0.339|RT @jeremyscahill: Trump's final tv ad is a masterpiece: https://t.co/DQK1ZIajP1
phiI94|twitter|0.6249|0.0|0.661|0.339|RT @jeremyscahill: Trump's final tv ad is a masterpiece: https://t.co/DQK1ZIajP1
divinetechinque|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
divinetechinque|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
AzadCandace|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
AzadCandace|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
OneTrump4All|joshgremillion|0.8745|0.0|0.63|0.37|RT @joshgremillion: Amazing support for @realDonaldTrump in NYC! Our driver is from Bangladesh and he is supporting Trump! #ElectionDay #MA
JakeLuciano1|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
JakeLuciano1|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
agentbar|BigT47119041|0.0|0.0|1.0|0.0|RT @BigT47119041: Donald Trump is putting it in your hands it all up you guys https://t.co/sB3QqKcrit
agentbar|twitter|0.0|0.0|1.0|0.0|RT @BigT47119041: Donald Trump is putting it in your hands it all up you guys https://t.co/sB3QqKcrit
SammieDolce|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
koogmo|emilysparkles|0.0|0.0|1.0|0.0|RT @emilysparkles: When an uneducated white dude literally invites shaming for voting for Trump on Facebook #GoHigh #ButSubtweetFirst https
mllsos7|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump now leading IN by 45 points.  RCP has him by 10.  Something is happening.
chrislewis_9|SirAbiola|0.0|0.0|1.0|0.0|RT @SirAbiola:  If Black People Voted For Donald Trump #ElectionDay https://t.co/QLqez43Rsv
chrislewis_9|amp|0.0|0.0|1.0|0.0|RT @SirAbiola:  If Black People Voted For Donald Trump #ElectionDay https://t.co/QLqez43Rsv
aussiedinos|doylething|0.0|0.0|1.0|0.0|RT @doylething: Some of the #ElectionNight games in London: Pussy Grabber and Trump Tower Jenga https://t.co/LdZWQRIJIc
aussiedinos|twitter|0.0|0.0|1.0|0.0|RT @doylething: Some of the #ElectionNight games in London: Pussy Grabber and Trump Tower Jenga https://t.co/LdZWQRIJIc
lisahatchet|johnlegend|0.0|0.0|1.0|0.0|"RT @johnlegend: Donald Trump is unfit for the office of president. Fortunately, there's an exceptionally qualified candidate @HillaryClinto"
bronxhenchmen|BonnieMadden|0.0|0.0|1.0|0.0|"RT @BonnieMadden: Once a crook, always a crook. VOTE TRUMP!"
HitchDied|JYSexton|-0.6874|0.294|0.706|0.0|"RT @JYSexton: If Trump freaks out and destroys the Trump Cake, this whole thing still wasn't worth it but..."
JocyTorralba|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
JocyTorralba|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
KiingMarc0|BrendanWHoward|0.5719|0.0|0.764|0.236|RT @BrendanWHoward: If trump wins I'll give $100 to 1 person who retweets this
Rub_Her_Toe|genesisbarzallo|0.6369|0.0|0.634|0.366|RT @genesisbarzallo: if you voted for trump please unfollow me thanks
_llisaaaa|tropicocunt|0.0|0.0|1.0|0.0|RT @tropicocunt: She voted for trump https://t.co/65kGJojFIv
_llisaaaa|twitter|0.0|0.0|1.0|0.0|RT @tropicocunt: She voted for trump https://t.co/65kGJojFIv
racfink47|jamessmurray|0.3802|0.08|0.747|0.172|Screw Donald Trump and Hillary Clinton! @jamessmurray definitely has my vote cuz I believe in him
parisscarlett94|trillmarn|-0.5994|0.178|0.822|0.0|@trillmarn soo what do you think trump or clinton who was pro war in iraq will do with presidency
Phillygr8|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
rcsummerall|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
TRINITYPRAISE|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
justwaldrop|WalshFreedom|-0.7876|0.338|0.558|0.104|"RT @WalshFreedom: I'm not saying this ELECTION is rigged, but Trump is right: The SYSTEM is rigged. Rigged to help Elites and rigged to s"
Makuna_4|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
TheRebelDelgado|br_uk|0.4767|0.0|0.763|0.237|RT @br_uk: Frank Lampard is fascinated by Donald Trump #ElectionDay https://t.co/ob4yyjAfPd
TheRebelDelgado|twitter|0.4767|0.0|0.763|0.237|RT @br_uk: Frank Lampard is fascinated by Donald Trump #ElectionDay https://t.co/ob4yyjAfPd
errrmaryam|Lord_Sugar|0.0|0.0|1.0|0.0|"RT @Lord_Sugar: can be @piersmorgan assistant in the executive loos at the white house. Piers hands Trump toilet roll, Nigel wipes https://"
errrmaryam||0.0|0.0|1.0|0.0|"RT @Lord_Sugar: can be @piersmorgan assistant in the executive loos at the white house. Piers hands Trump toilet roll, Nigel wipes https://"
swinshi|voxdotcom|0.3818|0.0|0.874|0.126|RT @voxdotcom: There are five people alive who have ever been president. None of them voted for Trump. https://t.co/7nufIhy28Y
swinshi|vox|0.3818|0.0|0.874|0.126|RT @voxdotcom: There are five people alive who have ever been president. None of them voted for Trump. https://t.co/7nufIhy28Y
ericvtine|ironghazi|0.5859|0.0|0.833|0.167|RT @ironghazi: Wow. Venn diagram showing Trump Voters (blue) and People Who Have Said The N Word This Week (yellow) https://t.co/amaQ9l8qzK
ericvtine|twitter|0.5859|0.0|0.833|0.167|RT @ironghazi: Wow. Venn diagram showing Trump Voters (blue) and People Who Have Said The N Word This Week (yellow) https://t.co/amaQ9l8qzK
Fatfufu_|nbc4i|0.0|0.0|1.0|0.0|RT @nbc4i: 102-year-old woman casts her vote for Donald Trump. https://t.co/rhJNJSy0rf https://t.co/jmz9hMN9YY
Fatfufu_|nbc4i|0.0|0.0|1.0|0.0|RT @nbc4i: 102-year-old woman casts her vote for Donald Trump. https://t.co/rhJNJSy0rf https://t.co/jmz9hMN9YY
InvestmentClubB|conservativetribune|0.7579|0.0|0.606|0.394|Hours Before Polls Close Supreme Court Gives Trump MASSIVE Good News https://t.co/a2IMrXT7DA
dalton_arfman98|saintpiercing|0.0|0.0|1.0|0.0|RT @saintpiercing: Retweet if you'd rather this pickle be president than Donald Trump https://t.co/PYVVwYBpXN
dalton_arfman98|twitter|0.0|0.0|1.0|0.0|RT @saintpiercing: Retweet if you'd rather this pickle be president than Donald Trump https://t.co/PYVVwYBpXN
Reckless__Alex|GavinFree|0.128|0.0|0.941|0.059|RT @GavinFree: I've been waiting to wake up from a dream for months now but I don't think it's going to happen. This trump thing is totally
DarrenjMcLaren|BritishVogue|0.0|0.0|1.0|0.0|RT @BritishVogue: The US Election: What Happens When? https://t.co/sD7EYjbzX3 #ElectionDay https://t.co/ofAJuyfF1k
DarrenjMcLaren|vogue|0.0|0.0|1.0|0.0|RT @BritishVogue: The US Election: What Happens When? https://t.co/sD7EYjbzX3 #ElectionDay https://t.co/ofAJuyfF1k
vampedexo|trapsouIed|0.5719|0.0|0.821|0.179|RT @trapsouIed: If Trump   Wins The Election I Am Moving   Out Of The Country  Goodbye   America   Hello   EXO PLANET
piercebboop|TheDonaldNews|0.627|0.0|0.708|0.292|RT @TheDonaldNews: LOOK AT CURRENT POPULAR VOTE!! TRUMP ==&gt;&gt; 6600  HILLARY===&gt;2043
laurie6805|rnlisa64|0.0|0.0|1.0|0.0|RT @rnlisa64: Voted Trump!!! #MAGA https://t.co/FTWASnfuRJ
laurie6805|twitter|0.0|0.0|1.0|0.0|RT @rnlisa64: Voted Trump!!! #MAGA https://t.co/FTWASnfuRJ
Margojs|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
cvrlosflores|YG|-0.5719|0.371|0.479|0.15|"RT @YG: All trump supports unfollow me, &amp; Suck my dick"
ariewestahl_2|WORLDSTAR|0.8126|0.0|0.519|0.481|RT @WORLDSTAR: If Trump wins vs. If Hilary wins https://t.co/pjJmaLZJjI
ariewestahl_2|twitter|0.8126|0.0|0.519|0.481|RT @WORLDSTAR: If Trump wins vs. If Hilary wins https://t.co/pjJmaLZJjI
MillyOdlum|EwanGreenwood|0.7351|0.0|0.78|0.22|RT @EwanGreenwood: Jokes that out of 350 million+ people in the US literally the best they could come up with was Trump and Clinton
Brisxyda|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
Brisxyda|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
bubblezhangpop|scamfuI|0.4404|0.0|0.775|0.225|@scamfuI imagine how many trump supporters will get in your mentions
olimpiadazayts1|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
olimpiadazayts1|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
SON_DJunior|TracyFortShow|0.636|0.0|0.811|0.189|"RT @TracyFortShow: I loved when Mr. Khan said, ""Mr. Trump this is not YOUR America, this is OUR America!'. https://t.co/EJg8bWLayb"
SON_DJunior|twitter|0.636|0.0|0.811|0.189|"RT @TracyFortShow: I loved when Mr. Khan said, ""Mr. Trump this is not YOUR America, this is OUR America!'. https://t.co/EJg8bWLayb"
Donwood72|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Donald #Trump. Follow @nbcconnecticut for the latest election news.https://t.co/zFdT7UCG1F
_WesleyRose|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
_WesleyRose|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
mtnbvan|davidcommon|-0.9417|0.515|0.485|0.0|@davidcommon @CBCGloria Horrible. And why letting Trump continually incite such violence &amp; harassment has been so irresponsible. Predictable
MadddieA19|caitlyngalinac_|0.7469|0.085|0.637|0.278|"RT @caitlyngalinac_: Idc if you like trump or clinton, but I have no respect for you if you call ppl that like a candidate you don't ""stupi"
mytq1354|erwoti|0.5622|0.0|0.752|0.248|RT @erwoti: Who is BETTER for the world?Vote and RT Widely#ElectionDay#voted#myvote2016#ElectionNight #WTFAmericaIn5WordsTrump
ALANDexter2020|MattGertz|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
ALANDexter2020|twitter|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
haugherin|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
Avionn2|BettyFckinWhite|0.0|0.0|1.0|0.0|"RT @BettyFckinWhite: By the way, if Trump gets elected, nothing you can do, folks. Although the Hitler Time Travel people, maybe there is."
GJoelChury|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
TrumpDyke|CROWENATION2016|0.4374|0.0|0.874|0.126|RT @CROWENATION2016: Calling all MILITARY in Pensacola!  Trump needs #FL panhandle to rise! Please contact everyone &amp; tell them to get
shalyseea|spkhp|0.0772|0.0|0.947|0.053|RT @spkhp: Me: who are you voting forKinder: TrumpMe: whyKinder: because he wants to send me back to Africa and I want to goMe: https:/
shalyseea||0.0772|0.0|0.947|0.053|RT @spkhp: Me: who are you voting forKinder: TrumpMe: whyKinder: because he wants to send me back to Africa and I want to goMe: https:/
CNC_Tethis|MattGertz|-0.7054|0.295|0.705|0.0|@MattGertz Tapper is an idiot. The whole of CNN can't be trusted. Trump doesn't lie either.
MiRobinette|troyesivan|-0.3182|0.133|0.867|0.0|RT @troyesivan: i dont mean to be a tease but....like...imagine not having to hear about donald trump anymore 
LibraChronicles|libertytarian|-0.6486|0.238|0.762|0.0|"RT @libertytarian: Seriously, even though Janet Reno died yesterday,I wonder who she's voting for todayDemocrat in Florida after all@Re"
Ayethatsmera|CjayyTaughtHer|0.0|0.0|1.0|0.0|RT @CjayyTaughtHer: Trump Vs Hillary  https://t.co/e3XUMJbgFY
Ayethatsmera|twitter|0.0|0.0|1.0|0.0|RT @CjayyTaughtHer: Trump Vs Hillary  https://t.co/e3XUMJbgFY
faketrentford|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
soph2124|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
DR_DRE_a|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
sleepybaekhyun|twitter|0.0|0.0|1.0|0.0|my dad out here wearing his 'i voted' sticker after voting for trump https://t.co/pLPUbeFAZQ
ThomasAHester2|spkhp|-0.3724|0.164|0.836|0.0|RT @spkhp: Me: what do you know about TrumpKinder: Donald Trump doesn't respect women
ermagerdcamila|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
TroyConway10|twitter|0.0|0.0|1.0|0.0|TRUMP!! https://t.co/tsRNxln6R4
UJournalism|EmilyMiller|0.4574|0.0|0.857|0.143|RT @EmilyMiller: I'll be live on @OANN all #ElectionNight from Trump NYC party. Tune in for the latest! https://t.co/umIpjVDrjO
UJournalism|twitter|0.4574|0.0|0.857|0.143|RT @EmilyMiller: I'll be live on @OANN all #ElectionNight from Trump NYC party. Tune in for the latest! https://t.co/umIpjVDrjO
elaineolsen|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
PattyCamps2|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
mcwhirter81|LilDwat|0.6774|0.0|0.626|0.374|RT @LilDwat: @DebAlwaystrump trump is winning but don't stop voting! That's what they want!
britasticuk|MartinShkreli|0.5719|0.0|0.829|0.171|"RT @MartinShkreli: If Trump wins, my entire unreleased music collection, including unheard Nirvana, Beatles, and of course, Wu-Tang, comes"
7bugglettes|kurteichenwald|0.4588|0.0|0.889|0.111|"RT @kurteichenwald: 43. In 2007, Trump said his favorite book was his own, The Art of the Deal. Once he started running 4 president, he sai"
sazonova_silva|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
sazonova_silva|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
INFOS_EN|aol|-0.4939|0.211|0.789|0.0|Nevada judge rejects Trump request for order over early voting - AOL News https://t.co/XMuXmylUND
FilipDobi|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump now leading IN by 45 points.  RCP has him by 10.  Something is happening.
_ellietripp|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
Paulhardingjr|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: 90% of America does not approve of Congress &amp; Washington DC. Trump will DRAIN THE SWAMP! #MAGA
KidJaxn|twitter|-0.5423|0.171|0.829|0.0|"trump said he'll go back to the ""black fountain &amp; white fountain"" fuck it i'm out #ElectionNight https://t.co/s6CFeBSrHp"
Stevelubbesmey1|realalexjones|0.2263|0.0|0.863|0.137|Video: Machine Refuses to Allow Vote For Trump in Pennsylvania https://t.co/fPEIVXkkVg via @realalexjones
Stevelubbesmey1|infowars|0.2263|0.0|0.863|0.137|Video: Machine Refuses to Allow Vote For Trump in Pennsylvania https://t.co/fPEIVXkkVg via @realalexjones
MoodyliciousSpa|rweingarten|0.4404|0.0|0.868|0.132|RT @rweingarten: Must read @ezraklein: Donald Trumps candidacy is the first time American politics has left me truly afraid https://t.co/3
MoodyliciousSpa|twitter|0.4404|0.0|0.868|0.132|RT @rweingarten: Must read @ezraklein: Donald Trumps candidacy is the first time American politics has left me truly afraid https://t.co/3
FOX5Atlanta|fox5atlanta|0.0|0.0|1.0|0.0|Former President George W. Bush didn't vote for Trump or Clinton https://t.co/BkoURf2iqP #YouDecideFOX5 #FOX5atl
andrialisa24|chrislhayes|-0.5256|0.159|0.841|0.0|RT @chrislhayes: Trump is already laying the groundwork to contest the legitimacy of the election and it's incredibly dangerous.
jrwsjs|recordonline|0.1027|0.112|0.759|0.129|RT @recordonline: Trump spent a good portion of Election Day sowing doubt about the legitimacy of the election results https://t.co/zdp7B41
jrwsjs|t|0.1027|0.112|0.759|0.129|RT @recordonline: Trump spent a good portion of Election Day sowing doubt about the legitimacy of the election results https://t.co/zdp7B41
vmetu|YoungDems4Trump|-0.2244|0.178|0.618|0.204|RT @YoungDems4Trump: Lol the DNC just called me to see if I voted I said hell yeah I voted... for DONALD J TRUMP!#MAGA
mindoflauren|twitter|0.1139|0.0|0.88|0.12|i'm not sorry in saying you should not vote for trump because you will be sorry if you do https://t.co/dNo0IPTXH5
ChilesMedios|NaomiAKlein|-0.5707|0.228|0.685|0.087|RT @NaomiAKlein: 1 reason to crush #Trump? The climate crisis. I made this film w/ @GuardianAus abt whats at stake. Please watch! https://
ChilesMedios||-0.5707|0.228|0.685|0.087|RT @NaomiAKlein: 1 reason to crush #Trump? The climate crisis. I made this film w/ @GuardianAus abt whats at stake. Please watch! https://
ASAPFurgal|Johnny_Blaz3|-0.7003|0.407|0.593|0.0|RT @Johnny_Blaz3: Latinos for Trump = Blacks for Slavery
4fathers4life|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
4fathers4life|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
therealdelariva|youtube|0.7345|0.0|0.531|0.469| I can't with these Trump supporters haha #StraightDumb #grabembythepussy ! https://t.co/Xzj2b6ODnJ
JudyCorradi|megynkelly|0.0|0.0|1.0|0.0|"RT @megynkelly: 18 electoral votes are up for grabs in #Ohio, and the states own Republican Gov. John Kasich says he did not vote for #Tru"
CobyBethea|KeithOlbermann|0.4019|0.219|0.365|0.416|@KeithOlbermann pretty awful. Just like the real Trump
anajelllyy|flawedfacade|0.0|0.0|1.0|0.0|RT @flawedfacade: Y'all talmbout a Trump presidency turning the clock back 500 years when in reality it'll turn the clock back less than 50
tangopublishing|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
tangopublishing|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
junecrotty|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump now leading IN by 45 points.  RCP has him by 10.  Something is happening.
Fayrraah|WeLoveRobDyrdek|0.4404|0.0|0.791|0.209|RT @WeLoveRobDyrdek: Jon Stewart and Donald Trump beef is funny af https://t.co/j1HsilMOlH
Fayrraah|twitter|0.4404|0.0|0.791|0.209|RT @WeLoveRobDyrdek: Jon Stewart and Donald Trump beef is funny af https://t.co/j1HsilMOlH
flanders292|MSNBC|0.34|0.125|0.625|0.25|@MSNBC that video just proves that Trump supporters are stupid Hit the number button as the clear directions say to do
AnonBruja|voxdotcom|-0.7003|0.293|0.707|0.0|RT @voxdotcom: A Nevada judge gave the Trump campaigns voter fraud paranoia the smackdown it deserved https://t.co/AVCo4Dtjkl
AnonBruja|vox|-0.7003|0.293|0.707|0.0|RT @voxdotcom: A Nevada judge gave the Trump campaigns voter fraud paranoia the smackdown it deserved https://t.co/AVCo4Dtjkl
Cam_Cheetah|ImToBlame|0.8503|0.0|0.571|0.429|"RT @ImToBlame: ""OMG TRUMP WON KENTUCKY??!!"" Yes nigga. Have you been to Kentucky?"
AdrianConradie|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
AdrianConradie|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
len_volkel|shootist2015|0.0|0.0|1.0|0.0|"RT @shootist2015: #Trump smashing #CrookedHillary in early exit poll data from Naples, FL https://t.co/WfaoP82jYN"
len_volkel|naplesnews|0.0|0.0|1.0|0.0|"RT @shootist2015: #Trump smashing #CrookedHillary in early exit poll data from Naples, FL https://t.co/WfaoP82jYN"
Peraltafqw|ml|0.3182|0.134|0.63|0.236|Don't take life to seriously :) #nyvotes Hillary o Trump https://t.co/NTS4bGxIpA
Diggydou|youtube|0.3612|0.0|0.857|0.143|T is for TrumpGravity lets the chips fall where they may just like Dominoeffect. https://t.co/UfY4bEVaCp via @youtube
Diggydou|youtube|0.3612|0.0|0.857|0.143|T is for TrumpGravity lets the chips fall where they may just like Dominoeffect. https://t.co/UfY4bEVaCp via @youtube
_sadsquatch|revlfrixnds|0.3612|0.143|0.606|0.251|RT @revlfrixnds: the fact that trump actually has a chance to win makes me sick to my stomach
Jthemovielover|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
_lorenaax3|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
_lorenaax3|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
princessnnaay|Gloful_|-0.6486|0.301|0.699|0.0|RT @Gloful_: If you voted for Donald trump ya moms a whore
philmonaco67|LindaSuhler|0.6776|0.0|0.798|0.202|"RT @LindaSuhler: Your SINGLE VOTE could be the difference between Donald J. Trump winning or not.Whatever it takes, VOTE!!!!#VoteTrump"
phyllisinirmo|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
wilycyotee|twitter|0.0772|0.0|0.944|0.056|I just want to know what they would have done if their wives didn't voted for Trump? Aren't votes supposed to be pr https://t.co/Nc5V7dnnTc
scorpiotiger77|MarkUrban01|-0.0258|0.212|0.579|0.208|"RT @MarkUrban01: Yes indeed - and Trump's campaign manager has just retaliated, blaming republican establishment for lack of support #Elect"
echoezofsilence|jaureologist|-0.0516|0.207|0.591|0.202|RT @jaureologist: I DON'T CARE HOW MUCH Y'ALL HATE BOTH CANDIDATES YOU WILL VOTE FOR HILLARY WHETHER YOU LIKE IT OR NOT I REFUSE TO LET TRU
BrianRodd6|RealPika|0.4926|0.0|0.79|0.21|RT @RealPika: Pikachu would be better than Donald Trump and Hillary Clinton! https://t.co/Q5ZdbSHID2
BrianRodd6|twitter|0.4926|0.0|0.79|0.21|RT @RealPika: Pikachu would be better than Donald Trump and Hillary Clinton! https://t.co/Q5ZdbSHID2
yaboifortemps|Suxting|-0.2023|0.306|0.463|0.231|RT @Suxting: Dress up like a slutty Trump.
TerrynRob|DiamondandSilk|0.0|0.0|1.0|0.0|"RT @DiamondandSilk: There's only one man who wants to totally work for and put the American people first, that man is @realDonaldTrump. Vo"
tekusaaleksand2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
tekusaaleksand2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
LoredoLeslie|SheHatesJacoby|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
LoredoLeslie|twitter|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
nataweejunks|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
hmay26|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
hmay26|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
pmcg|TeaPainUSA|0.0|0.0|1.0|0.0|"RT @TeaPainUSA: Remember how just Kellyanne Conway called Trump's campaign an ""Act of Charity?""  Beer's cheaper at Yankee stadium.  https:/"
pmcg||0.0|0.0|1.0|0.0|"RT @TeaPainUSA: Remember how just Kellyanne Conway called Trump's campaign an ""Act of Charity?""  Beer's cheaper at Yankee stadium.  https:/"
__300___|J_valdebenito26|0.5719|0.0|0.837|0.163|RT @J_valdebenito26: If Trump wins I AM* a citizen so if you don't wanna get deported hmu so we can get married
TwittHappens|guinnesssud|0.3182|0.0|0.881|0.119|"@guinnesssud  Trump /O Keefe/ Obannon philosophy  2% truth, 98% misdirection and hyperbole.  Then tell as loud and https://t.co/Dm3VXKHqTo"
TwittHappens|twitter|0.3182|0.0|0.881|0.119|"@guinnesssud  Trump /O Keefe/ Obannon philosophy  2% truth, 98% misdirection and hyperbole.  Then tell as loud and https://t.co/Dm3VXKHqTo"
polishedoffinc|alaskantexanQCT|0.0|0.0|1.0|0.0|RT @alaskantexanQCT: Yo fam heading to Philly with some homies and 2 vans. Gonna take Black Trump voters 2 the polls ALL DAY tomorrow! #MAG
SamElizabethan|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
SamElizabethan|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
MarissaJo225|twitter|0.5719|0.0|0.448|0.552|If Trump* wins https://t.co/FarPb6q8l0
jillianmallory|Latina|0.743|0.102|0.59|0.308|"RT @Latina: ""It would be sweet, sweet justice if after every attack...it was the Latino vote that defeated Donald Trump."" -@ananavarro on @"
DLPaxt|DiamondandSilk|0.0|0.0|1.0|0.0|"RT @DiamondandSilk: .@realDonaldTrump is Americans only Choice.  Blacks, whites, Hispanics, Asian, Latinos  Vote, Vote, Vote. ......Vote Tr"
brittykittyj|brooklyn_alexa|0.0|0.0|1.0|0.0|RT @brooklyn_alexa: @TheGinger_KING trump 2016
brownryan6|JaredWyand|0.5859|0.128|0.667|0.206|RT @JaredWyand: It's simple...Trump needs NHIf he loses FL he needs PA &amp; MIIf he wins FL loses NC he needs MI or PAIf he wins FL he
mcloughh|TaraMeehan62|0.3612|0.0|0.737|0.263|RT @TaraMeehan62: Donald trump look like a fat carrot
flaw3d_b3auty|younggwhite|0.0|0.0|1.0|0.0|RT @younggwhite: imagine back in 08' if Obama had done even .0001 of what's surfaced about Trump. they would've burned him at the stake
MarthaDepuy|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
MarthaDepuy|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
TheGiantHogweed|clmazin|-0.8442|0.302|0.698|0.0|"RT @clmazin: ""Fail Bigly"" (2031) - Barry Pepper stars as failed Republican nominee Donald J. Trump in the story of his historic loss to Hil"
Biu1231|FrankLuntz|-0.5423|0.137|0.863|0.0|RT @FrankLuntz: The turnout in Madison and Ann Arbor suggest that Trump is going to have a bad time in Wisconsin and Michigan.  #ElectionNi
buffriku98|Astrofyre|-0.3612|0.238|0.762|0.0|RT @Astrofyre: RT for Arin ignore for Trump https://t.co/1vlI0SGuI2
buffriku98|twitter|-0.3612|0.238|0.762|0.0|RT @Astrofyre: RT for Arin ignore for Trump https://t.co/1vlI0SGuI2
YOCUMILA|chanddlerriggs|0.0|0.0|1.0|0.0|RT @chanddlerriggs: boys at my school: feminists are so triggered over everything lolme: i would rather have hillary than trumpboys at
BlazinHope|StarbucksSanae|0.2146|0.378|0.291|0.33|"@StarbucksSanae NO, DON'T LET TRUMP WIN, NO, DON'T LET HILLARY WIN! WE'RE SCREWED!"
ImALegendKiller|dormgod|0.5859|0.0|0.745|0.255|"RT @dormgod: Per the BBC, 17% excited about a Clinton presidency. 13% excited about a Trump presidency. #ElectionNight"
keating_eleanor|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
siqqest|Possum_Jones|-0.25|0.083|0.917|0.0|@Possum_Jones @sabbytappy I think you're alone on this one if you think trump has any prior knowledge of global politics. Nor do you itseems
kimulleuer|Joannahausmann|0.2732|0.0|0.884|0.116|RT @Joannahausmann: Neighbor: Who you vote for?Me: ClintonNeighbor: Well I'm voting Trump because Im an AmericanMe:....#ElectionDay htt
masahiko_x|Prince_Sakamaki|0.0|0.0|1.0|0.0|RT @Prince_Sakamaki: Kino is gayBut not for Trump 
DeeAlumni|BoxingHype|0.0|0.0|1.0|0.0|RT @BoxingHype: VIDEO: Conor McGregor goes off at Donald Trump.. #UFC205 https://t.co/GszVpWGz2a
DeeAlumni|twitter|0.0|0.0|1.0|0.0|RT @BoxingHype: VIDEO: Conor McGregor goes off at Donald Trump.. #UFC205 https://t.co/GszVpWGz2a
RockieBilbrey|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
RockieBilbrey|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
cristhianne28|jamesmichael|-0.2732|0.084|0.916|0.0|RT @jamesmichael: s/o to this golden moment where Trump let us all know that he doubted his own wife would vote for him. https://t.co/rDdUt
cristhianne28|t|-0.2732|0.084|0.916|0.0|RT @jamesmichael: s/o to this golden moment where Trump let us all know that he doubted his own wife would vote for him. https://t.co/rDdUt
icufromhere|DonaldJTrumpJr|0.5696|0.0|0.872|0.128|"RT @DonaldJTrumpJr: If you have friends in MI, OH, FL, PA -- CALL THEM and tell them to VOTE TRUMP! You can make a difference! #MAGA #Tru"
_nicholasgreen_|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
_nicholasgreen_|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
rabcyr|fronxer|0.4939|0.18|0.506|0.313|RT @fronxer: white men: well at least a trump win would be interesting hahahaliterally everybody else: no pls we're going to suffer and d
bob_smite|PunkDuck_|0.5719|0.0|0.709|0.291|RT @PunkDuck_: If Trump wins I'll upload ''How To Mercury''
deniza_gureva|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
deniza_gureva|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
tia6sc|trfgrp|0.0|0.0|1.0|0.0|"RT @trfgrp: Our projection: Trump 306 Clinton 223 w/CO, VA &amp; WI possibly breaking Trump as ""hidden voter"" #trumptiderolls https://t.co/u34D"
tia6sc|t|0.0|0.0|1.0|0.0|"RT @trfgrp: Our projection: Trump 306 Clinton 223 w/CO, VA &amp; WI possibly breaking Trump as ""hidden voter"" #trumptiderolls https://t.co/u34D"
vmwabe|YoungDems4Trump|-0.2244|0.178|0.618|0.204|RT @YoungDems4Trump: Lol the DNC just called me to see if I voted I said hell yeah I voted... for DONALD J TRUMP!#MAGA
ketch169|seangentille|-0.2714|0.211|0.635|0.154|"RT @seangentille: Thanks to Bill Belichick, you can hate the Patriots again! https://t.co/NlgtjTiwsM https://t.co/vtRDzNeEbf"
ketch169|sportingnews|-0.2714|0.211|0.635|0.154|"RT @seangentille: Thanks to Bill Belichick, you can hate the Patriots again! https://t.co/NlgtjTiwsM https://t.co/vtRDzNeEbf"
ranpaq|Cory_1077|0.0|0.0|1.0|0.0|RT @Cory_1077: VOTE TRUMP To get rid if the #PoliticalCorruption in our Country #MakeAmericaGreatAgain   #MakeAmer
purmetheus|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
terrydvl|szeachmoment|0.0772|0.0|0.885|0.115|RT @szeachmoment: @theglobaluniter @DonaldJTrumpJr panhandle dweller here. Everyone I know voted Trump.
dcfriend3|twitter|0.0|0.0|1.0|0.0|Boohoo-wait until president Trump starts investigating Hillary and all the others mentioned in the #wikileaks relea https://t.co/sBjizsa0kZ
AdamKeyes23|SheriffClarke|0.3612|0.0|0.706|0.294|@SheriffClarke praying your way to a Trump victory?
MariannBenway|ChristieC733|0.743|0.0|0.687|0.313|"RT @ChristieC733: Whatever you can do, I would appreciate. I say pray for me, I pray for you.""~ Donald Trump #ElectionFinalThoughts #G"
orendax|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
orendax|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
LySaundraJanee|twitter|0.6369|0.09|0.631|0.279|"It feels like ""Hunger Games Could Legitimately Be In Our Future If Donald Trump Wins"" Day https://t.co/Amy7Hicbqn"
MentalJargon|FatalAn0xia|0.0|0.0|1.0|0.0|"@FatalAn0xia Trump will be leading for ages, Red states close polls early as conservatives vote earlier in the day."
factiod|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
lamaramironova4|cosmopolitan|-0.0772|0.204|0.612|0.184|Trolls Attacked Trump's Website and the Results Are Hilarious https://t.co/ktIHc4CTNE https://t.co/1CldjekfdW
backwaterdogs|mitchellvii|0.34|0.0|0.893|0.107|"RT @mitchellvii: I expect Trump to win KY and IN, but not by 50 points.  We'll see if anything near that holds."
andurilprime|PeterSlattery3|0.0|0.0|1.0|0.0|"RT @PeterSlattery3: For a brief moment tonight, someone figured out that you could make Trump's website say... anything you wanted: https:/"
andurilprime||0.0|0.0|1.0|0.0|"RT @PeterSlattery3: For a brief moment tonight, someone figured out that you could make Trump's website say... anything you wanted: https:/"
punk_perkins|kylekinane|-0.2732|0.237|0.529|0.234|"RT @kylekinane: ""No matter what, get out and VOTE.""""Cool. I might go with a third party candidate/Trump.""""OH GOD DONT VOTE YOU'LL RUIN"
Kjslom5|AdelleNaz|0.0|0.0|1.0|0.0|"RT @AdelleNaz: Star-Spangled Banner being sung by diverse group of Americans in front of #HiltonMidtown, where Trump-Pence ElectionNight pa"
QGS24|EthanQuinn4|-0.1147|0.155|0.722|0.123|"RT @EthanQuinn4: Trump certainly isn't great, but just look at this. https://t.co/tfakDBWgg0"
QGS24|twitter|-0.1147|0.155|0.722|0.123|"RT @EthanQuinn4: Trump certainly isn't great, but just look at this. https://t.co/tfakDBWgg0"
alpha_joe86|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
ollgsheeran|ium44k|-0.5423|0.212|0.788|0.0|RT @ium44k: @screamgreys jovens que gravaram mil snaps falando fuck you trump me add
hotelco226|Dianne09314822|0.6093|0.0|0.834|0.166|"RT @Dianne09314822: Drove my 85 &amp; 90 year old friends to vote today!  Been married 65 years, they voted Trump!! https://t.co/x1kvjuHgmC"
hotelco226|twitter|0.6093|0.0|0.834|0.166|"RT @Dianne09314822: Drove my 85 &amp; 90 year old friends to vote today!  Been married 65 years, they voted Trump!! https://t.co/x1kvjuHgmC"
stevemeredith21|mitchellvii|0.5719|0.0|0.829|0.171|"RT @mitchellvii: Trump now up 23,000 including Indies in Pinellas County, FL.  In 2012, Obama won this by 26,000."
00LovelyDay00|vivelafra|0.0|0.0|1.0|0.0|RT @vivelafra: ATTENTION #TRUMPTRAIN: The MSM narrative is beginning to CRUMBLE.  States long given to #Hillary are now back in the toss-up
meganderson01|toriking68|0.7845|0.0|0.717|0.283|RT @toriking68: Everyone bashes Trump like Hillary is any better and everyone bashes Hillary like Trump is any better...in the end we're al
jaque_bauer|t|-0.1027|0.223|0.567|0.21|https://t.co/Rb06T0bEkPTHE RAG NAMED THE DAILY MAIL IS NOT FIT FOR USE AS FISH PAPER. ITS CLEARLY A COMMUNIST RAG OF  PROPAGANDA AND SHIT
ero_Ashley|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
ero_Ashley|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
OBauby|MsAmyHerron|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
OBauby|theguardian|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
wise_diva|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
wise_diva|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
JayySoWavyy|whoissizzIe|0.0|0.0|1.0|0.0|RT @whoissizzIe: This right here: Trump vs Clinton  https://t.co/Lzf7ghjFWY
JayySoWavyy|twitter|0.0|0.0|1.0|0.0|RT @whoissizzIe: This right here: Trump vs Clinton  https://t.co/Lzf7ghjFWY
SadMarchand|dril|0.0|0.0|1.0|0.0|RT @dril: if you ask me this election could end about 100 different ways:1) trump gets 0% of the vote2) trump gets 1% of the vote3) trum
krazyjake313|DiamondandSilk|0.0|0.0|1.0|0.0|"RT @DiamondandSilk: .@realDonaldTrump is Americans only Choice.  Blacks, whites, Hispanics, Asian, Latinos  Vote, Vote, Vote. ......Vote Tr"
Moratayaa61|DonDziesinski|0.0|0.066|0.868|0.066|RT @DonDziesinski: I feel like Trump &amp; Hilary are two divorced parents fighting over custody of us but we kinda just wanna go live with gra
Designertype|ananavarro|-0.2732|0.087|0.913|0.0|"RT @ananavarro: Hey Nevadans, u know why Trump is suing? To keep Hispanics from polls b/c he knows we're voting against him. Redouble your"
LoverofAll777|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
LoverofAll777|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
kristinrocksu2|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
kristinrocksu2|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
keepcalmila|TheFactsOfShade|-0.0516|0.216|0.588|0.196|RT @TheFactsOfShade: Donald Trump has no chance. https://t.co/Zl9lLtgFgT
keepcalmila|twitter|-0.0516|0.216|0.588|0.196|RT @TheFactsOfShade: Donald Trump has no chance. https://t.co/Zl9lLtgFgT
taylor_kayh|twitter|0.0|0.0|1.0|0.0|I meant she's (Judge) on to the Trump ppl asking for names.  Never give them names. https://t.co/kCiw8MDKWk
FaithAndorf|LeafyIsHere|0.4238|0.139|0.589|0.272|"RT @LeafyIsHere: If Trump wins I'll release nudes, not a joke"
PrisonUK|deray|-0.5106|0.125|0.875|0.0|"RT @deray: The @NYTimes has printed a list of all of the people, places, &amp; things that Trump has insulted on Twitter during the campaign. h"
rvacts|Jvmzie|0.0|0.0|1.0|0.0|"RT @Jvmzie: I'm going to bed. When I wake up, Donald Trump will be prime minister of America. You heard it here first people, I'm never wro"
coolinit81|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
coolinit81|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
VetCapitalist|JBellSATX|0.0|0.0|1.0|0.0|@JBellSATX @KGBVeteran @FrankLuntz Trump 282
randomsubu|twitter|0.0|0.0|1.0|0.0|"America to Trump, soon enough. https://t.co/juGgZWDt01"
Blondeadroit|oliverdarcy|0.5267|0.0|0.841|0.159|RT @oliverdarcy: Trump winning big in this Fox exit poll category: Can candidate bring change? *Clinton: 13%*Trump: 82% https://t.co/e1u
Blondeadroit|t|0.5267|0.0|0.841|0.159|RT @oliverdarcy: Trump winning big in this Fox exit poll category: Can candidate bring change? *Clinton: 13%*Trump: 82% https://t.co/e1u
JakeLuciano1|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
dkarnold|pittsburgh|0.0|0.0|1.0|0.0|Voting Issues: Some Trump Voters Reporting Ballots Switching To Clinton https://t.co/Akzyjb2cQ3
SylvieBommel|nytimes|0.5859|0.0|0.787|0.213|"The 1,024 Ways Clinton or Trump Can Win the Election - The New York Times https://t.co/Ake05mmtu6"
VSStangl|FrankLuntz|-0.5423|0.137|0.863|0.0|RT @FrankLuntz: The turnout in Madison and Ann Arbor suggest that Trump is going to have a bad time in Wisconsin and Michigan.  #ElectionNi
Zander9899|mimimayesTN|0.4019|0.0|0.863|0.137|@mimimayesTN @rharrisonfries @Reince @GOP collected millions in Trump's name ~ spent 0 to help Trump~Letter asking for donation from Reince
HalfABlueeSkyy|jamesmichael|-0.2732|0.084|0.916|0.0|RT @jamesmichael: s/o to this golden moment where Trump let us all know that he doubted his own wife would vote for him. https://t.co/rDdUt
HalfABlueeSkyy|t|-0.2732|0.084|0.916|0.0|RT @jamesmichael: s/o to this golden moment where Trump let us all know that he doubted his own wife would vote for him. https://t.co/rDdUt
starsabove0oru|flawedfacade|0.0|0.0|1.0|0.0|RT @flawedfacade: Y'all talmbout a Trump presidency turning the clock back 500 years when in reality it'll turn the clock back less than 50
MoweryRoger|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
laraherrick|someecards|0.0|0.0|1.0|0.0|RT @someecards: Trump mixed up 'county' and 'country' on the day he could be elected to run one of those things. https://t.co/ThAsXQXKlx ht
laraherrick|someecards|0.0|0.0|1.0|0.0|RT @someecards: Trump mixed up 'county' and 'country' on the day he could be elected to run one of those things. https://t.co/ThAsXQXKlx ht
raymarin96|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
raymarin96|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
61Rinaldi|hockeydeb21|-0.4466|0.257|0.616|0.128|RT @hockeydeb21: LEAKED CLINTON INTERNAL DOCUMENT: Discourage Trump Supporters with Bogus Polls and Declaring Election Over https://t.co/cJ
61Rinaldi|t|-0.4466|0.257|0.616|0.128|RT @hockeydeb21: LEAKED CLINTON INTERNAL DOCUMENT: Discourage Trump Supporters with Bogus Polls and Declaring Election Over https://t.co/cJ
WilliamSDraper|JRehling|-0.3612|0.116|0.884|0.0|RT @JRehling: Donald Trump started life with a $14 million loan from his father.He thinks the system is rigged against him.#ElectionNight
gravenoise|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
jBSTEEL_|ironghazi|0.5859|0.0|0.833|0.167|RT @ironghazi: Wow. Venn diagram showing Trump Voters (blue) and People Who Have Said The N Word This Week (yellow) https://t.co/amaQ9l8qzK
jBSTEEL_|twitter|0.5859|0.0|0.833|0.167|RT @ironghazi: Wow. Venn diagram showing Trump Voters (blue) and People Who Have Said The N Word This Week (yellow) https://t.co/amaQ9l8qzK
jg1935|breitbart|0.8016|0.0|0.675|0.325|Pat Caddell on Whatever It Takes: Trump Wins Because The People Want Their Country Back https://t.co/gWSLqTFkrW I hope Caddell is right!
HHAWKBOSS|America_1st_|0.3578|0.0|0.829|0.171|RT @America_1st_: BREAKINGMachine Refuses to Allow Vote For Trump in Pennsylvania!!#VoterFraud #ElectionDay https://t.co/f5efnGdWF3
HHAWKBOSS|twitter|0.3578|0.0|0.829|0.171|RT @America_1st_: BREAKINGMachine Refuses to Allow Vote For Trump in Pennsylvania!!#VoterFraud #ElectionDay https://t.co/f5efnGdWF3
HandToForehead|WendyBrandes|0.0|0.0|1.0|0.0|@WendyBrandes  Trump brought Melania here illegally as a sex slave.
Pam55561059|megynkelly|0.2023|0.0|0.921|0.079|"RT @megynkelly: .@marthamaccallum: In terms of top the quality for a candidate, change is very impt to voters tonight. 82% of voters are g"
radronin|twitter|0.7627|0.0|0.432|0.568|C'mon guys support Trump! Support America!!! https://t.co/smj92ECnHE
ashkeylim|Mcbrownie|0.3612|0.0|0.906|0.094|"RT @Mcbrownie: Texas had a wave of crickets, it's been raining for like a week strait, Trump is leading in some polls, ITS THE END OF TIMES"
feoktistkondra7|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
feoktistkondra7|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
wtfstavo|ladygaga|0.5106|0.0|0.87|0.13|RT @ladygaga: Emma from Wisconsin has Cerebral Palsy. In a wheelchair her whole life. She saw the video of Trump making fun of a disabled r
luckydbldd|mrbeercrusher|0.0|0.0|1.0|0.0|RT @mrbeercrusher: Expect a Trump victory in North Carolina announced around eight o'clock eastern time. Trump up 3.7% in the average of ex
alex__dalton96|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
alex__dalton96|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
JesslcaHansen_|Hope012015|0.3818|0.0|0.898|0.102|"RT @Hope012015: Kellyanne Conway just said on msnbc that Trump will accept the results tonight, ""As he sees them,"" she wouldn't say what th"
wells1780|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
OliviaArntzen|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
awoll2016|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
CurlsGawd|Y2SHAF|0.6597|0.076|0.694|0.229|RT @Y2SHAF: If Donald Trump wins the presidency with no background in politics I shouldn't have to graduate university to get a good job in
tmoroney4697|WhySharksMatter|0.6124|0.0|0.773|0.227|"RT @WhySharksMatter: I was just informed that Jews should forgive anti-Semitic Trump supporters because ""it's the Christian thing to do""."
Xamerican|MariaYes2trump|0.81|0.108|0.514|0.378|RT @MariaYes2trump: TRUMP VOTER LINES ARE HUGE! THERE IS NO WAY HILLARY CAN LEGALLY WIN! https://t.co/ImNnufMQAi via @wordpressdotcom
Xamerican|themarshallreport|0.81|0.108|0.514|0.378|RT @MariaYes2trump: TRUMP VOTER LINES ARE HUGE! THERE IS NO WAY HILLARY CAN LEGALLY WIN! https://t.co/ImNnufMQAi via @wordpressdotcom
Dirtyassbum|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
Dirtyassbum|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
m_abagail|NBCNews|0.296|0.098|0.758|0.144|RT @NBCNews: Can Trump pull an upset in Virginia? The state has been a key to every GOP president's win since 1924: https://t.co/F2MLlKpC7Y
m_abagail|nbcnews|0.296|0.098|0.758|0.144|RT @NBCNews: Can Trump pull an upset in Virginia? The state has been a key to every GOP president's win since 1924: https://t.co/F2MLlKpC7Y
standupkid|costareports|0.0|0.0|1.0|0.0|"RT @costareports: On the phone w/ Giuliani. He just left Trump's apt. Said Trump is ""watching everything even tho I'm telling him not to."""
_gigi_vega|TheMexicanVines|0.6597|0.0|0.795|0.205|"RT @TheMexicanVines: If you voted for Trump today, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why th"
zeabraa|polaroidbones|-0.607|0.184|0.816|0.0|RT @polaroidbones: DONT SPLIT THE DEMOCRATIC VOTE TOMORROW CAUSE YOU DONT WANNA BE STUCK HILLARY OR TRUMP! ITS ONLY GONNA LEAVE US WITH TRU
adelaidakirill3|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
adelaidakirill3|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
lukey1223|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
GirlCountry33|politicususa|0.3182|0.0|0.892|0.108|RT @politicususa: Caught on Camera: Donald Trump Makes Sure His Own Wife Votes For Him via @politicususa https://t.co/3kCNKprMMX #p2 #ctl
GirlCountry33|politicususa|0.3182|0.0|0.892|0.108|RT @politicususa: Caught on Camera: Donald Trump Makes Sure His Own Wife Votes For Him via @politicususa https://t.co/3kCNKprMMX #p2 #ctl
maxxbadazzent|GLOGangHQ|0.0|0.0|1.0|0.0|RT @GLOGangHQ: Donald Trump Hillary Clinton Chief Keef GO VOTE TODAY CHIEF KEEF 4 PRESIDENT #Election2016 #MyVote2016 https://t.co/
maxxbadazzent|t|0.0|0.0|1.0|0.0|RT @GLOGangHQ: Donald Trump Hillary Clinton Chief Keef GO VOTE TODAY CHIEF KEEF 4 PRESIDENT #Election2016 #MyVote2016 https://t.co/
NatetheBRD|brianstelter|0.0|0.0|1.0|0.0|"RT @brianstelter: Lara Trump just confirmed on @CNN that ""Melania and I both voted for Donald Trump"" https://t.co/hHaCkCVsjX"
NatetheBRD|twitter|0.0|0.0|1.0|0.0|"RT @brianstelter: Lara Trump just confirmed on @CNN that ""Melania and I both voted for Donald Trump"" https://t.co/hHaCkCVsjX"
Brad4rdHay|onlxn|0.3041|0.0|0.899|0.101|RT @onlxn: CONWAY: What's with the cake?TRUMP: Little tradition I have. I like to mark big life events by eating Rutger Hauer https://t.co
Brad4rdHay|t|0.3041|0.0|0.899|0.101|RT @onlxn: CONWAY: What's with the cake?TRUMP: Little tradition I have. I like to mark big life events by eating Rutger Hauer https://t.co
Neto_Bruck|Enrique_Acevedo|0.0|0.0|1.0|0.0|RT @Enrique_Acevedo: Trump finally got his wall. #TheLatinoVote
Lofdaproduction|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Lofdaproduction|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
CoppedNews|washingtonpost|-0.5859|0.241|0.759|0.0|"#coppednews The Fix: Donald Trump's Election Day insinuations of voter fraud, explained https://t.co/DeLPwh74PL"
GenineU|DonaldJTrumpJr|0.4939|0.0|0.849|0.151|RT @DonaldJTrumpJr: Independent and late breaking voters heading towards Trump. Our voters are inspired to take back America. Incredible. P
OlavPonomaryov|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
OlavPonomaryov|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ts65136|TheTrumpLady|0.3786|0.095|0.754|0.151|"RT @TheTrumpLady: #Trump LOOKIN' GOOD Already! Wait for the WORKING CLASS, NEW VOTERS, &amp; 15% UNDECIDED To Come Home &amp; Vote! #TrumpTrain #Tr"
peachymarz|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
theylovehannah_|flawedfacade|0.0|0.0|1.0|0.0|RT @flawedfacade: Y'all talmbout a Trump presidency turning the clock back 500 years when in reality it'll turn the clock back less than 50
yoonirim|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
selinakrieg|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Hail_Tisa|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Hail_Tisa|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
patchrhythm|thecreatorgee|0.5267|0.0|0.702|0.298|RT @thecreatorgee: i can't believe trump is winning inna south
jscandiffwow|thehill|-0.5358|0.308|0.692|0.0|"RT @thehill: Tom Brady's wife: No, we don't support Trump https://t.co/bpcKrcVzXL https://t.co/rcYriClzgz"
jscandiffwow|thehill|-0.5358|0.308|0.692|0.0|"RT @thehill: Tom Brady's wife: No, we don't support Trump https://t.co/bpcKrcVzXL https://t.co/rcYriClzgz"
QopperP|twitchytrex|-0.3541|0.193|0.657|0.149|"RT @twitchytrex: legit im so worried about women, poc, and lgbt+ rights if Trump wins all the shit ive seen with mike pence makes me want t"
aydooon|FNLOPPC|0.4019|0.091|0.705|0.203|RT @FNLOPPC: Know that Hilary and Trump have no power. The true Power is in the hands of God. #GodIsThere
thanroberts|DaRealDanBaulch|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
thanroberts|t|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
biebsdemz|David16996|-0.4215|0.167|0.833|0.0|RT @David16996: How can people defend trump after all his comments about women ugh  #ElectionNight
beccaw__|champagneomar|0.6597|0.0|0.722|0.278|RT @champagneomar: All these Trump supporters look like they would be the first ones to purge
CesarMonroyO|YouTube|0.4753|0.0|0.781|0.219|I liked a @YouTube video from @thunderf00t https://t.co/eMJvHdFUo1 Trump vs Clinton: The FINAL showdown!
CesarMonroyO|youtube|0.4753|0.0|0.781|0.219|I liked a @YouTube video from @thunderf00t https://t.co/eMJvHdFUo1 Trump vs Clinton: The FINAL showdown!
theyloveflacko|Imskeno|-0.2617|0.311|0.444|0.244|"RT @Imskeno: Trump trash, but he funny as shit"
MG_LilChris|_Latishhaaaa|-0.5423|0.243|0.757|0.0|RT @_Latishhaaaa: I'm just gonna leave this right here .. Trump is such an idiot  https://t.co/Qd0G85Znt2
MG_LilChris|twitter|-0.5423|0.243|0.757|0.0|RT @_Latishhaaaa: I'm just gonna leave this right here .. Trump is such an idiot  https://t.co/Qd0G85Znt2
ra_estella|religiouscaviar|0.743|0.0|0.751|0.249|"RT @religiouscaviar: Hillary's been serving looks since the 60s, and tonight she'll serve Trump and his supporters by winning the presidenc"
calvalais|ProgtopiaBooks|0.0|0.0|1.0|0.0|RT @ProgtopiaBooks: Some Pittsburgh machines changing from Trump to Hillary.Problems call 1-866-OUR-VOTE
ovchinn78750209|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ovchinn78750209|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
Tommy_Reason|twitter|0.5719|0.0|0.654|0.346|Me if Trump wins:Me if Hillary wins: https://t.co/jbKJp1LaBw
MichaelMcGan|VickiMDonovan|-0.8155|0.361|0.639|0.0|"RT @VickiMDonovan: #california Pay NO attention to exit polls, they're FAKE, designed to keep you from voting TRUMP!"
AllenAdkins2|LindaSuhler|0.6776|0.0|0.798|0.202|"RT @LindaSuhler: Your SINGLE VOTE could be the difference between Donald J. Trump winning or not.Whatever it takes, VOTE!!!!#VoteTrump"
aubraleigh|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
aubraleigh|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
BurovaLyutseya|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
BurovaLyutseya|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
notbapecamo|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
notbapecamo|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
sofiadaviddd|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
CoxaleeLee|mitchellvii|0.5859|0.0|0.759|0.241|RT @mitchellvii: Pat Caddell: I think Trump will win todays voting by a large margin.https://t.co/zqJNzOaS2m
purplestar2015|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump will get between 35 and 40% of the Hispanic vote.
jennyy882|memeprovider|-0.1695|0.196|0.804|0.0|"RT @memeprovider: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
ChristineIs43|bakedalaska|0.4225|0.16|0.621|0.219|RT @bakedalaska: I am so proud to have voted for Donald J. Trump today. Couldn't be happier. Thank you everyone for your support. #MAGASe
H93Chris|CarltonBarrass|0.3612|0.0|0.884|0.116|RT @CarltonBarrass: 'Choosing between trump or clintons like choosing either jerry or kate mccann to watch the bairns for u'
BrexitAftermath|MightyBusterBro|0.0|0.0|1.0|0.0|RT @MightyBusterBro: .A MUST SEE VIDEOINSPIRATIONAL MOMENTFINAL TRUMP RALLY@realDonaldTrump#VOTE  #ElectionDay #MyVote2016 #MAGA htt
kendallbrown491|ViraI|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
kendallbrown491|twitter|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
_nataliaduran|Enrigr8|-0.4588|0.115|0.885|0.0|RT @Enrigr8: If u in the 20% of Latinos that voted for Trump u are hereby banned from eating pernil or dancing salsa/bachata ever again htt
catovitch|nihilistwaraxe|0.0|0.0|1.0|0.0|"@nihilistwaraxe Trump will make them use qwerty, finally"
nataliyamaksim7|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
nataliyamaksim7|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
maryzimnik|GuardianUS.|0.6369|0.0|0.792|0.208|Best place to get the #returns: @GuardianUS. Follow live #Election2016 updates as #votes come in | #ImWithHer    https://t.co/gJ2xFimRPK
maryzimnik|theguardian|0.6369|0.0|0.792|0.208|Best place to get the #returns: @GuardianUS. Follow live #Election2016 updates as #votes come in | #ImWithHer    https://t.co/gJ2xFimRPK
pmswolfy|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
chrisldoster|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
joeycongi98|twitter|-0.1531|0.15|0.726|0.124|Don't try and tell me that Clinton is a good Candidate. Just as bad as Trump in my opinion. https://t.co/qZ1mmkSkjQ
USA_with_Trump|docdhj|0.0|0.0|1.0|0.0|RT @docdhj: I have lived in Michigan for 32 years &amp; have never seen the lines as long as today! A Sea of Red! @realDonaldTrump @AJDelgado13
JR777771|LeslieMarshall|0.0|0.0|1.0|0.0|RT @LeslieMarshall: It's official! #DonaldTrump has made history!  https://t.co/ijA6W9utx5.#TaxReturns #ImWithHer #NeverTrump #ElectionDay
JR777771|t|0.0|0.0|1.0|0.0|RT @LeslieMarshall: It's official! #DonaldTrump has made history!  https://t.co/ijA6W9utx5.#TaxReturns #ImWithHer #NeverTrump #ElectionDay
ayu_lestari128|FaZeZubZer|-0.4019|0.316|0.526|0.158|RT @FaZeZubZer: Idk why people support Donald trump he is racist. #ElectionNight
Vadersleash|speechboy71|-0.5106|0.202|0.798|0.0|RT @speechboy71: If only Trump had insulted the spouses of every Republican #whatcouldhavebeen https://t.co/ElY8QxJL3U
Vadersleash|twitter|-0.5106|0.202|0.798|0.0|RT @speechboy71: If only Trump had insulted the spouses of every Republican #whatcouldhavebeen https://t.co/ElY8QxJL3U
SamsonovNodar|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
SamsonovNodar|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
BidiBidiDemDem|GRlFFERS|-0.3612|0.244|0.565|0.191|"RT @GRlFFERS: This Trump Supporter just turned around and told me ""have fun in conversion therapy fag"" wtf omg https://t.co/klMNKR9l8e"
BidiBidiDemDem|twitter|-0.3612|0.244|0.565|0.191|"RT @GRlFFERS: This Trump Supporter just turned around and told me ""have fun in conversion therapy fag"" wtf omg https://t.co/klMNKR9l8e"
cpopa2001|thetigersez|0.3612|0.0|0.889|0.111|RT @thetigersez: Donald Trump's face always looks like a toddler's who has just pooped in the potty for the first time. https://t.co/oZMqG9
cpopa2001|t|0.3612|0.0|0.889|0.111|RT @thetigersez: Donald Trump's face always looks like a toddler's who has just pooped in the potty for the first time. https://t.co/oZMqG9
ManuelTunzer_|twitter|0.6908|0.0|0.659|0.341|Green&amp;socialist party 6% #trump 7% #clinton 63% bei #electionparty in #vienna :) https://t.co/MnRBLSZ88j
MattM3502|RawStory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
MattM3502|rawstory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
DrBenWhitham|dmuleicester|0.0|0.0|1.0|0.0|RT @dmuleicester: #ElectionDay: DMU expert predicts the first 100 days for Trump &amp; Clinton: https://t.co/e8Zo6qWhYr https://t.co/2pRMHGA1kH
DrBenWhitham|dmu|0.0|0.0|1.0|0.0|RT @dmuleicester: #ElectionDay: DMU expert predicts the first 100 days for Trump &amp; Clinton: https://t.co/e8Zo6qWhYr https://t.co/2pRMHGA1kH
speccymcspec|OwensDamien|-0.561|0.256|0.646|0.099|"RT @OwensDamien: Lets hope the closing shot of this terrible movie is Trump all alone in his gold apartment, realising hes forgotten his"
_ogluis1|bIakout|0.0|0.0|1.0|0.0|RT @bIakout: The White House if Trump becomes President. https://t.co/2ekd9vwLlr
_ogluis1|twitter|0.0|0.0|1.0|0.0|RT @bIakout: The White House if Trump becomes President. https://t.co/2ekd9vwLlr
MRileygautier|ZachingOff_|-0.5423|0.283|0.594|0.123|RT @ZachingOff_: If you think people who support Trump are racists you're part of the problem
mswilliams1|TMZ|-0.69|0.343|0.592|0.065|RT @TMZ: Donald Trump Tower Barricaded By Dump Trucks To Prevent Attacks! https://t.co/1fCw13uwgq
mswilliams1|twitter|-0.69|0.343|0.592|0.065|RT @TMZ: Donald Trump Tower Barricaded By Dump Trucks To Prevent Attacks! https://t.co/1fCw13uwgq
aNickel4thought|dyfl|0.0|0.0|1.0|0.0|"RT @dyfl: Just when you think this election cannot possibly offer up any more gifts to the meme economy, here comes Cake Trump"
JoSheram|jerome_corsi|-0.5859|0.153|0.847|0.0|RT @jerome_corsi: TRUMP NEEDS ALL POSSIBLE VOTERS IN PA - voter fraud being reported EVENING HOURS WILL DECIDE ELECTION - get all Trump vot
lionsboi|twitter|-0.6419|0.243|0.673|0.084|"Trump is a vile person with a litany of flaws to numerous to mention. Cory is just a prick, I wouldn't piss on him https://t.co/CXDw9ntFcR"
anthonytaylor_|eddyrivas|0.5927|0.0|0.862|0.138|"RT @eddyrivas: I try not to do this too much on social media, but I will say I hope we never hear from Donald Trump in a political setting"
sadmexicanchica|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
mags_holes|dubstep4dads|0.0|0.0|1.0|0.0|RT @dubstep4dads: trump: what are you drawingmelania: uhh... nothing https://t.co/2EMzgUx8yc
mags_holes|twitter|0.0|0.0|1.0|0.0|RT @dubstep4dads: trump: what are you drawingmelania: uhh... nothing https://t.co/2EMzgUx8yc
_Timone|ClarenceJWhite|0.0|0.069|0.863|0.069|RT @ClarenceJWhite: I feel like Trump &amp; Hillary are two divorced parents fighting over custody of us but we kinda just wanna go live with g
MitchellA_12|JaredWyand|0.1511|0.0|0.935|0.065|RT @JaredWyand: Donald Trump #voted in NYC!5 rallies yesterday and the man was up at 6am doing shows. I want a worker in the White House.
AG_Conservative|twitter|-0.3612|0.186|0.688|0.126|"Again, Trump now only guaranteed ""amnesty,"" but also made border security unpopular. He hurt every cause he claimed https://t.co/STvWBNLTmZ"
trade420|Thomas1774Paine|-0.3612|0.122|0.878|0.0|RT @Thomas1774Paine: #Trump Voters Complain Their Votes Locked Out of Electronic Voting Machines in New York **RT**RT**RT** #voterfraud htt
AlissaLeighh_|__ImNotReal__|0.1779|0.088|0.797|0.116|RT @__ImNotReal__: No we're voting against trump cause he's a despicable human being. If we had a better option than Hillary we'd vote agai
Indiiaaa15|polaroidbones|-0.607|0.184|0.816|0.0|RT @polaroidbones: DONT SPLIT THE DEMOCRATIC VOTE TOMORROW CAUSE YOU DONT WANNA BE STUCK HILLARY OR TRUMP! ITS ONLY GONNA LEAVE US WITH TRU
TimGriffin02061|costareports|0.3612|0.0|0.848|0.152|@costareports even Trump doesn't listen to Rudy. See Trump is like the rest of us
CathySalmons|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
grahamfthoran|BornToWin____|0.0|0.0|1.0|0.0|RT @BornToWin____: So Trump Jr came to speak at my school today and this was the results https://t.co/7GhiRC9Ryl
grahamfthoran|twitter|0.0|0.0|1.0|0.0|RT @BornToWin____: So Trump Jr came to speak at my school today and this was the results https://t.co/7GhiRC9Ryl
Saya_relativity|hstcaahs|-0.9381|0.463|0.495|0.042|RT @hstcaahs: @Hope012015 @latimes trump will go to his grave lying! He just can't help himself! Just never stops lying! Crooked Lying #dru
pdowdski|Queen_Caleb|-0.1761|0.115|0.8|0.084|RT @Queen_Caleb: The fact that straight people really don't see that big of a deal of a Trump/Pence presidency...Y'all really lack empath
Cmoneymontana|RonnieFieg|0.5719|0.0|0.764|0.236|"RT @RonnieFieg: If Trump wins, going to relocate the team to Kith Canada."
essar1|FrankConniff|-0.4767|0.134|0.866|0.0|RT @FrankConniff: Trump campaign crying foul over reports that flagrant acts of democracy are happening in precincts all over the country.
minikennirusso|tillery_13|0.7003|0.0|0.691|0.309|RT @tillery_13: I support Trump and I have just as many black friends as I do white https://t.co/UeQpCygEqL
minikennirusso|twitter|0.7003|0.0|0.691|0.309|RT @tillery_13: I support Trump and I have just as many black friends as I do white https://t.co/UeQpCygEqL
kevhazel33|foxandfriends|0.5927|0.0|0.806|0.194|"RT @foxandfriends: .@GovMikeHuckabee: Hillary Clinton needs celebrities to get a crowd, but Donald Trump's supporters aren't coming for a f"
HannahHoelzen|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
myhorsecowboy|RichardGrenell|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
myhorsecowboy|twitter|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
EloyChronicles|MailOnline|-0.6124|0.238|0.762|0.0|"Some much needed distraction from a long and tense ballot counting night. Trump in a robe, anyone?  https://t.co/eaeOd3Ywhr via @MailOnline"
EloyChronicles|dailymail|-0.6124|0.238|0.762|0.0|"Some much needed distraction from a long and tense ballot counting night. Trump in a robe, anyone?  https://t.co/eaeOd3Ywhr via @MailOnline"
coldplayitcool|jaureologist|-0.0516|0.207|0.591|0.202|RT @jaureologist: I DON'T CARE HOW MUCH Y'ALL HATE BOTH CANDIDATES YOU WILL VOTE FOR HILLARY WHETHER YOU LIKE IT OR NOT I REFUSE TO LET TRU
_Uncreative_16|__Chona__|0.1531|0.092|0.764|0.143|"RT @__Chona__: Everyone has the right to vote for who they want. Getting tired of the ""if it was your friend you wouldn't let them vote for"
dericdunk|DRUDGE_REPORT|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: PA VOTERS REPORT SEEING TRUMP VOTES SWITCH TO CLINTON BEFORE THEIR EYES... https://t.co/ZSKfysoxkE
dericdunk|pittsburgh|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: PA VOTERS REPORT SEEING TRUMP VOTES SWITCH TO CLINTON BEFORE THEIR EYES... https://t.co/ZSKfysoxkE
ragwed12|JOMainEvent|0.7081|0.0|0.754|0.246|"RT @JOMainEvent: I don't know about you guys, but this is crucial! We all know Trump supporters want Change!#ElectionNight #voted #TeamT"
PantsuitEnFuego|JMilesColeman|0.0|0.0|1.0|0.0|"RT @JMilesColeman: Floyd County, where KY House Speaker Stumbo (D) hails from, is going 70% Trump. Was 54% Conway in #KYGov. #kyelect #kyvo"
ocstangmanck|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
Rub_Her_Toe|SuperDuperHunt|0.0|0.0|1.0|0.0|RT @SuperDuperHunt: Me when I first heard Trump was running vs. me today #ElectionDay https://t.co/anv5MSLik9
Rub_Her_Toe|twitter|0.0|0.0|1.0|0.0|RT @SuperDuperHunt: Me when I first heard Trump was running vs. me today #ElectionDay https://t.co/anv5MSLik9
LinWeeks|LilDwat|0.6774|0.0|0.626|0.374|RT @LilDwat: @DebAlwaystrump trump is winning but don't stop voting! That's what they want!
davebucknut|LindaSuhler|0.0|0.0|1.0|0.0|"RT @LindaSuhler: TUESDAY, NOV 08, 2016DONALD J. TRUMP VICTORY PARTYDonald J. Trump &amp; Governor Mike Pence7 PM ET New York, NYhttps://t.c"
Peinert16|Sporf|-0.3182|0.173|0.827|0.0|RT @Sporf: BREAKING: Stone Cold interrupts the Donald Trump rally.  #ElectionDay( @thrillis4)https://t.co/zJZAmoHlNY
Peinert16|twitter|-0.3182|0.173|0.827|0.0|RT @Sporf: BREAKING: Stone Cold interrupts the Donald Trump rally.  #ElectionDay( @thrillis4)https://t.co/zJZAmoHlNY
Odangles|bbydev_|-0.5859|0.272|0.625|0.103|"@bbydev_ trump is for sure giant douche, clinton is turd sandwich because shes always full of shit"
c6ron|youtube|-0.3237|0.152|0.848|0.0|OMG! JAMES COMEY WONT SLEEP TONIGHT AFTER WHAT TRUMP JUST EXPOSED ABOUT HIM https://t.co/zojhHga1oA
RyzaJem|boomitsmaia|-0.34|0.362|0.638|0.0|RT @boomitsmaia: i swear trump has no political background?
librtytakngroot|varepall|0.7824|0.0|0.735|0.265|RT @varepall: OHIO IS LOOKING GOOD FR TRUMP.  THANK YOU OHIO FOR GETTING OUT THE VOTES.  KEEP THEM COMING.POLLS ARE OPEN
PennyLDuncan|WDFx2EU8|0.0|0.0|1.0|0.0|"RT @WDFx2EU8: THIS FUCKING WHITE, HETEROSEXUAL, COLLEGE-EDUCATED, LIBERAL-ARTS MAJOR FROM ILLINOIS JUST VOTED FOR TRUMP! MAGA!!!!!!!!!! #IV"
aalyanxkhan|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
aalyanxkhan|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
kiamarie30|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
tonimcen|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Medievalgirltoo|SandyWarf|-0.4019|0.119|0.881|0.0|RT @SandyWarf: I SMELL #Trump Victory in the air  If  you encounter any problems voting #ElectionDay call VOTER ASSISTANCE HOTLINE to re
SadeJKing|TheFamilyAlpha|-0.1779|0.131|0.764|0.105|"RT @TheFamilyAlpha: Things are looking good for Trump, regardless of the outcome of this race, The Family Alpha will continue to provide po"
blvckpyrvmxd|hokagemaria|-0.2732|0.255|0.576|0.169|RT @hokagemaria: Donald trump did a great job exposing the racism that we are constantly told doesn't exist.
PGongola|jko417|0.0|0.0|1.0|0.0|"RT @jko417: ""Donald Trump is not the person that the media has depicted him to be"" #Trump2016 (Vine by @USAforTrump2016) https://t.co/R3G7K"
PGongola|t|0.0|0.0|1.0|0.0|"RT @jko417: ""Donald Trump is not the person that the media has depicted him to be"" #Trump2016 (Vine by @USAforTrump2016) https://t.co/R3G7K"
96Wille|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
96Wille|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
jeanne_tall|0hour|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
jeanne_tall|twitter|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
mattelmonsoon|nxswitch|0.5719|0.0|0.619|0.381|RT @nxswitch: me if trump wins https://t.co/QEXkf8UI8V
mattelmonsoon|twitter|0.5719|0.0|0.619|0.381|RT @nxswitch: me if trump wins https://t.co/QEXkf8UI8V
kristinaswaffo1|PriceParker2|-0.8126|0.346|0.654|0.0|"RT @PriceParker2: If voting for Trump makes you a racist, does voting for Hillary make you a criminal?"
ariatriplex|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
ariatriplex|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Matoozie|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
Matoozie|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
dmoore564|larrymeath|-0.0276|0.093|0.818|0.089|RT @larrymeath: It's difficult to sneer at a nation who may very well put #Trump in White House   when your own nation has Boris Johnson a
leoxva_|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
leoxva_|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
imwithh3r|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
imwithh3r|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
hakbooty|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
LeahR77|mitchellvii|0.5719|0.0|0.85|0.15|"RT @mitchellvii: Romney won Brevard County by 36,000 votes in 2012.  I calculate Trump leads it by 52,000 votes.  +16,000 votes for Trump o"
DearNormaa|cosmo_8a|0.0258|0.148|0.7|0.152|RT @cosmo_8a: If trump wins and anybody starts a riot let me know I'm trying to get a tv or something
illestclev|AweeBurrEee|-0.8594|0.263|0.737|0.0|RT @AweeBurrEee: people who oppose Hillary talk about her stance on abortion but won't discuss Trump's child rape case?????? babies are bab
Vazquez__Javier|LeafyIsHere|0.4238|0.139|0.589|0.272|"RT @LeafyIsHere: If Trump wins I'll release nudes, not a joke"
throughthatmist|ilysmarigrande|0.6393|0.076|0.7|0.224|"RT @ilysmarigrande: Hillary might not be the best candidate, but u can't deny that she's better than Trump. I urge you to vote tomorrow. #I"
mattleto1|NS_swiat|0.0|0.0|1.0|0.0|@NS_swiat have I said I wanted trump ? Try again
Shade58b|mitchellvii|0.4404|0.0|0.805|0.195|"RT @mitchellvii: Trump leads IND 72-25.  Good Lord people, something is happening here."
GrayDeenShaka|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
GrayDeenShaka|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
BruceMezistrano|RebellionReport|0.128|0.092|0.797|0.112|"RT @RebellionReport: If Trump loses, tell your kids after three SCOTUS appointments you satisfied their life and country for your self righ"
CarolPe91164590|thejoshuablog|0.0|0.0|1.0|0.0|RT @thejoshuablog: Voters For Trump Ad https://t.co/N9w4cHQcXg #BasketOfDeplorables
CarolPe91164590|youtube|0.0|0.0|1.0|0.0|RT @thejoshuablog: Voters For Trump Ad https://t.co/N9w4cHQcXg #BasketOfDeplorables
Toridevon|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
Toridevon|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
TJrasar|WaysThingsWork|0.1695|0.0|0.886|0.114|RT @WaysThingsWork: Obama endorsing Hillary and bashing trump? Let's not forget about this https://t.co/olDwdXaYFB
TJrasar|twitter|0.1695|0.0|0.886|0.114|RT @WaysThingsWork: Obama endorsing Hillary and bashing trump? Let's not forget about this https://t.co/olDwdXaYFB
tlvrp_russia|therussophile|-0.6908|0.322|0.678|0.0|"#Moscow #SaintPetersburg WikiLeaks criticizes both Hillary Clinton and Donald Trump, condemns McCarthyite Russia https://t.co/LWkUgemgl5"
gusmac2|1visionamd|0.0|0.0|1.0|0.0|RT @1visionamd: @nationdivided  many Democrats are voting for Trump to!
whomadewho102|RealVinnieJames|0.7213|0.0|0.768|0.232|RT @RealVinnieJames: TRUMP SUPPORTERS WHO HAVE NOT VOTED: Stay OUT of the Twitter trending column. That's where the head games are played.
switt1181|SemperFiCop|-0.7034|0.245|0.755|0.0|RT @SemperFiCop: #ImVotingBecause Donald Trump has been fighting for us against the corrupt establishment. TOMORROW WE FIGHT FOR HIM #Drain
c446591fcb1a479|juanitamoutlaw|0.0|0.0|1.0|0.0|RT @juanitamoutlaw: @DonaldJTrumpJr @JudyMichiganMomIM SAYIN IT LOUD!I VOTED @realDonaldTrump !AND I'M PROUD!NO Trump signs so I MADE M
sweatyglow|brujaaverde|-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
sweatyglow||-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
DawnSwe12515208|mitchellvii|0.7998|0.0|0.736|0.264|RT @mitchellvii: The last RCP Poll had Trump winning KY by 17.  He is currently winning by 52 points.Monster vote?  Dem crossovers?
krispy126|RickyRapsFL|0.0|0.0|1.0|0.0|RT @RickyRapsFL: RT if you voted for Donald J. Trump for president! #TrumpTheVote #ElectionDay #ElectionNight https://t.co/hlfCUbHHM8
krispy126|twitter|0.0|0.0|1.0|0.0|RT @RickyRapsFL: RT if you voted for Donald J. Trump for president! #TrumpTheVote #ElectionDay #ElectionNight https://t.co/hlfCUbHHM8
lastname_jeter|Kxngjorden|0.0|0.0|1.0|0.0|RT @Kxngjorden: Trump Trump Trump
PRsH0mbr3|SemperFiCop|-0.7034|0.245|0.755|0.0|RT @SemperFiCop: #ImVotingBecause Donald Trump has been fighting for us against the corrupt establishment. TOMORROW WE FIGHT FOR HIM #Drain
CindyCallinsky|Bill_Cimbrelo|0.8777|0.0|0.653|0.347|RT @Bill_Cimbrelo: @TweetingYarnie I voted Stein here. I know you went Trump. It's all good - anyone but a Clinton! Good luck to the USA an
akaMJz|PsyQo_Kolby|0.6249|0.0|0.541|0.459|@PsyQo_Kolby now I kinda want trump to fucking win 
Brendag38323989|Right_Smarts|0.0|0.0|1.0|0.0|RT @Right_Smarts: Scientific Poll Shows Trump With Yuge Lead in Swing States https://t.co/srwK0AEO5M #Trump2016
Brendag38323989|infowars|0.0|0.0|1.0|0.0|RT @Right_Smarts: Scientific Poll Shows Trump With Yuge Lead in Swing States https://t.co/srwK0AEO5M #Trump2016
KatieHedley69|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
KatieHedley69|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
espizzzzle|vPabIito|0.3182|0.176|0.543|0.281|RT @vPabIito: Yo when Trump wins I'm ready for this Civil War 2 I stay strapped https://t.co/sI6k9cUmrd
espizzzzle|twitter|0.3182|0.176|0.543|0.281|RT @vPabIito: Yo when Trump wins I'm ready for this Civil War 2 I stay strapped https://t.co/sI6k9cUmrd
JBDorward|dve1198|0.7845|0.0|0.603|0.397|RT @dve1198: Trusting Donald Trump with America is like trusting David Moyes with Man Utd
harrysuckszayn|pattonoswalt|0.0|0.0|1.0|0.0|RT @pattonoswalt: OMG Donald Trump just texted this to me. Does he already know I voted for Clinton? https://t.co/7COBWg7imR
harrysuckszayn|twitter|0.0|0.0|1.0|0.0|RT @pattonoswalt: OMG Donald Trump just texted this to me. Does he already know I voted for Clinton? https://t.co/7COBWg7imR
Robirdie23|Lexual__|-0.4588|0.143|0.857|0.0|"RT @Lexual__: Also, Trump has very shady business dealings that involved forced labor and discriminating against black tenants. Again.... B"
aznuman|GaryLineker|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
aznuman|twitter|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
ImMoonMan|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
ImMoonMan|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
holaitsangiexo|yvetteposts|0.0|0.0|1.0|0.0|RT @yvetteposts: for the 20% of the latinos voting for trump: ya moms a hoe https://t.co/SIsGBxji1L
holaitsangiexo|twitter|0.0|0.0|1.0|0.0|RT @yvetteposts: for the 20% of the latinos voting for trump: ya moms a hoe https://t.co/SIsGBxji1L
RadicalRW|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
mariizzle_|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
OZZWALD_1|SadderDre|0.5719|0.0|0.764|0.236|RT @SadderDre: if Trump wins I'll PayPal everyone a chicken wing that RTs this.
greatoneAKIRA|TheSuplexCity|0.0|0.0|1.0|0.0|RT @TheSuplexCity: Message to Donald Trump! https://t.co/nSd7K97SGa
greatoneAKIRA|twitter|0.0|0.0|1.0|0.0|RT @TheSuplexCity: Message to Donald Trump! https://t.co/nSd7K97SGa
Matriiix_RL|BrendanWHoward|0.5719|0.0|0.764|0.236|RT @BrendanWHoward: If trump wins I'll give $100 to 1 person who retweets this
Sports_Guy50|britishbullybee|0.5719|0.0|0.654|0.346|@britishbullybee I was saying that if trump wins ......
LowKiiiiSavage|YahBoyJiraiya|0.0|0.0|1.0|0.0|RT @YahBoyJiraiya: RT for the Pervy SageLike for Donald Trump  https://t.co/ZlznSSSkNm
LowKiiiiSavage|twitter|0.0|0.0|1.0|0.0|RT @YahBoyJiraiya: RT for the Pervy SageLike for Donald Trump  https://t.co/ZlznSSSkNm
StevensResa|carlajo1947|0.0|0.0|1.0|0.0|RT @carlajo1947: REPORTS ARE COMING OUT THAT MICHIGAN VOTING IS CURRENTLY A LANDSLIDE VICTORY FOR TRUMP! https://t.co/eFiVAidr9l
StevensResa|twitter|0.0|0.0|1.0|0.0|RT @carlajo1947: REPORTS ARE COMING OUT THAT MICHIGAN VOTING IS CURRENTLY A LANDSLIDE VICTORY FOR TRUMP! https://t.co/eFiVAidr9l
biyaf_A|facebook|0.0|0.0|1.0|0.0|Michelle Obama spent a lot of 2016 slaying Donald J. Trump without ever using his name https://t.co/DIkAqkmm34
HazelOsterhout|tpartynews|0.5411|0.0|0.857|0.143|"RT @tpartynews: Reince Priebus: Dont believe the garbage you read, were gonna put Trump in the White House &amp; save this country!""#Electi"
_evaax0|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_evaax0|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
hellohln|SoniaAnanti|0.0|0.0|1.0|0.0|RT @SoniaAnanti: Dont tell Trump: #Minnesota is about to elect a pioneering Somali-American Muslim woman https://t.co/ncKrRUiv35 #Election
hellohln|thenation|0.0|0.0|1.0|0.0|RT @SoniaAnanti: Dont tell Trump: #Minnesota is about to elect a pioneering Somali-American Muslim woman https://t.co/ncKrRUiv35 #Election
BJA1021|WeNeedTrump|0.25|0.0|0.857|0.143|RT @WeNeedTrump: Convince one more person today why we need Trump. #ElectionDay https://t.co/d8q3qpzVs3
BJA1021|twitter|0.25|0.0|0.857|0.143|RT @WeNeedTrump: Convince one more person today why we need Trump. #ElectionDay https://t.co/d8q3qpzVs3
in_myselff|PrisonPlanet|0.0258|0.14|0.679|0.181|"RT @PrisonPlanet: Reports out of Ohio at one polling station Trump supporters furious: Votes being flipped to Clinton, police called, allow"
ONLYTRUMP4USA|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
slmorris555|IankarloV16|0.4404|0.0|0.847|0.153|RT @IankarloV16: We Latinos are Family One Family Against Trump #imwithher #LoveTrumpsHate  #latinosvote thanks to all latinos
Spotdogs3|RickyRapsFL|0.0|0.0|1.0|0.0|RT @RickyRapsFL: RT if you voted for Donald J. Trump for president! #TrumpTheVote #ElectionDay #ElectionNight https://t.co/hlfCUbHHM8
Spotdogs3|twitter|0.0|0.0|1.0|0.0|RT @RickyRapsFL: RT if you voted for Donald J. Trump for president! #TrumpTheVote #ElectionDay #ElectionNight https://t.co/hlfCUbHHM8
blackwood_julie|DavidCornDC|-0.7096|0.312|0.688|0.0|RT @DavidCornDC: I have been banned by @realDonaldTrump. I was denied credentials for Trump election night event.
whiotv|Ohio_Politics|0.5719|0.0|0.778|0.222|RT @Ohio_Politics: .@HillaryClinton comments on what she'll do if she wins #ElectionNight https://t.co/9W2vgsBovh https://t.co/E7pUfLndti
whiotv|daytondailynews|0.5719|0.0|0.778|0.222|RT @Ohio_Politics: .@HillaryClinton comments on what she'll do if she wins #ElectionNight https://t.co/9W2vgsBovh https://t.co/E7pUfLndti
nimzaj_ruiz|drearetano|0.1371|0.102|0.741|0.157|RT @drearetano: for all of u voting for trump don't even  bother comin to invitational tryna score some tamales. tryna play my mom dirty li
daytondailynews|Ohio_Politics|0.5719|0.0|0.778|0.222|RT @Ohio_Politics: .@HillaryClinton comments on what she'll do if she wins #ElectionNight https://t.co/9W2vgsBovh https://t.co/E7pUfLndti
daytondailynews|daytondailynews|0.5719|0.0|0.778|0.222|RT @Ohio_Politics: .@HillaryClinton comments on what she'll do if she wins #ElectionNight https://t.co/9W2vgsBovh https://t.co/E7pUfLndti
rahcassi|LilTimye|0.0|0.0|1.0|0.0|RT @LilTimye: Whoever voted for trump ya moms a hoe
severianpolyak2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
severianpolyak2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
springfieldnews|Ohio_Politics|0.5719|0.0|0.778|0.222|RT @Ohio_Politics: .@HillaryClinton comments on what she'll do if she wins #ElectionNight https://t.co/9W2vgsBovh https://t.co/E7pUfLndti
springfieldnews|daytondailynews|0.5719|0.0|0.778|0.222|RT @Ohio_Politics: .@HillaryClinton comments on what she'll do if she wins #ElectionNight https://t.co/9W2vgsBovh https://t.co/E7pUfLndti
z1o9z6e9|NPR|0.0|0.0|1.0|0.0|RT @NPR: A spokesman for former President George W. Bush confirms to NPR that he and his wife voted for neither Donald Trump nor Hillary Cl
dasya_nesterova|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
dasya_nesterova|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
designdetails16|MeganSmiles|0.765|0.0|0.625|0.375|RT @MeganSmiles: Watch @LouDobbs on @FoxBusiness -much better &amp; he loves Trump  https://t.co/0muGdef3YZ
designdetails16|twitter|0.765|0.0|0.625|0.375|RT @MeganSmiles: Watch @LouDobbs on @FoxBusiness -much better &amp; he loves Trump  https://t.co/0muGdef3YZ
RealKidPoker|sawmillthug|0.4995|0.0|0.823|0.177|@sawmillthug they aren't deplorable. The ones who actually LIKE Trump are. 100% of them are deplorable.
Trillnfinesse|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
Trillnfinesse|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
papa_smurf34|SuspendedShaaa|0.9299|0.0|0.367|0.633|RT @SuspendedShaaa: @CNN Hilary will win or trump will win good luck !
smallant|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
smallant|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
r0ma_invicta|Thomas1774Paine|-0.3612|0.122|0.878|0.0|RT @Thomas1774Paine: #Trump Voters Complain Their Votes Locked Out of Electronic Voting Machines in New York **RT**RT**RT** #voterfraud htt
EledaReeth|rblandford|-0.5574|0.31|0.69|0.0|RT @rblandford: Shit. Sunderland South have gone for Trump.
RightAsRain7|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
RightAsRain7|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
trappinxc|ObamaSpotify|-0.5423|0.226|0.774|0.0|RT @ObamaSpotify: President Obama is currently listening to Fuck Donald Trump by YG
philmonaco67|surfermom77|-0.2263|0.101|0.899|0.0|RT @surfermom77: Undecided Voters 4 TrumpToday is the DAY we are going to take our country back &amp; #MakeAmericaGreatAgain#Vote4Trumphttps
impertinent78|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
impertinent78|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
alenaangel16|raaaqcity|0.5707|0.0|0.817|0.183|"RT @raaaqcity: please exercise your right to vote tomorrow! unless you're a trump supporter, then election day is on nov. 28th for you guys"
kenzdelrey|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
itistj1|twitter|0.7865|0.0|0.565|0.435|What Hillary will look like when she realizes TRUMP WON  https://t.co/td3SM5IFgt
beckypike34|farrightgregy|0.0|0.0|1.0|0.0|"RT @farrightgregy: RT RT_com: 1% reporting in - #Trump leading in early poll results in Kentucky, New Hampshire, Indiana #ElectionNig http"
naarwien|imskytrash|0.3089|0.0|0.852|0.148|RT @imskytrash: TRUMP: who are you voting forMELANIA: none of your damn business https://t.co/feCBRLKitX
naarwien|twitter|0.3089|0.0|0.852|0.148|RT @imskytrash: TRUMP: who are you voting forMELANIA: none of your damn business https://t.co/feCBRLKitX
TravisSeirer|DRUDGE_REPORT|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: PA VOTERS REPORT SEEING TRUMP VOTES SWITCH TO CLINTON BEFORE THEIR EYES... https://t.co/ZSKfysoxkE
TravisSeirer|pittsburgh|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: PA VOTERS REPORT SEEING TRUMP VOTES SWITCH TO CLINTON BEFORE THEIR EYES... https://t.co/ZSKfysoxkE
thgirtla|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
Kid_Codi_D|madirockssocks|0.7865|0.141|0.54|0.319|"@madirockssocks how hard would it have been to say ""hey trump I wish you the BEST of luck today"" tho? It's just unnecessary negativity."
ThaMoneyMonster|ABCDavidd|-0.5423|0.467|0.533|0.0|RT @ABCDavidd: Fuck Donald Trump
h8breeding|CherOfficiaI|0.6633|0.0|0.783|0.217|RT @CherOfficiaI: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
tam_raww|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
tam_raww|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
oxnfre|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
LaneMorrow10|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
LaneMorrow10|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
richardshadow1|AlysiaStern|-0.5553|0.146|0.854|0.0|"RT @AlysiaStern: @ananavarro My Hispanic family voted for TRUMP! You don't represent us, in fact you don't REPRESENT. Great work keeping yo"
DeplorableStorm|nationdivided|0.128|0.0|0.919|0.081|RT @nationdivided: Breaking news: Broward County Florida a democratic stronghold Republican turnout up 6% Democrat turnout down 6% that's a
zauxier|jimgeraghty|0.7351|0.0|0.714|0.286|"RT @jimgeraghty: The Trump party victory cake. This election is like a surreal, twisted dream where nothing makes sense and its taking f"
ThorntonMcEnery|twitter|0.0|0.0|1.0|0.0|"You guys, is Trump's concession going to be a Cirque du Soleil joint? https://t.co/6JJpJ0HlK2"
DCofStaff|LOLGOP|0.0516|0.138|0.714|0.148|RT @LOLGOP: EXIT POLL: 3 in 10 Trump supporters had trouble finding the exit to the polls.
panamahat1961|mitchellvii|0.3182|0.0|0.723|0.277|RT @mitchellvii: Trump leads Kentucky 77-20. :-)
thrashiva|JYSexton|-0.6874|0.294|0.706|0.0|"RT @JYSexton: If Trump freaks out and destroys the Trump Cake, this whole thing still wasn't worth it but..."
n_amaryllis|ViraI|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
n_amaryllis|twitter|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
thechubbstaa|abc15|-0.25|0.083|0.917|0.0|"RT @abc15: LIVE VIDEO: Protest at North High School -- students walked out to urge voters not to vote for Trump, Arpaio: https://t.co/OXDzd"
thechubbstaa|t|-0.25|0.083|0.917|0.0|"RT @abc15: LIVE VIDEO: Protest at North High School -- students walked out to urge voters not to vote for Trump, Arpaio: https://t.co/OXDzd"
_arivna|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
Saamprater|tpartynews|0.5411|0.0|0.857|0.143|"RT @tpartynews: Reince Priebus: Dont believe the garbage you read, were gonna put Trump in the White House &amp; save this country!""#Electi"
121536Mi|twitter|0.0|0.0|1.0|0.0|TheDebrief : 82% of Americans believe Donald Trump 'Can Bring Change'. But what sort of ch https://t.co/2xz0EZSHfZ) https://t.co/On3LQfweXI
Pudding_Brains_|GaryLineker|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
Pudding_Brains_|twitter|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
SheilaNJ|twitter|0.5927|0.109|0.64|0.25|OMG and this moron will have a job in the WH if Trump was to win. The man is already half senile. God help us all. https://t.co/tYatFgRMQZ
KopylovZoriy|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
KopylovZoriy|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
katkrchniak|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
LKGNanci|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
krazaykay_|TaylaaWayla_|-0.4404|0.23|0.599|0.17|RT @TaylaaWayla_: the fact that donald trump got a chance of winning goes to show ya tht america still white and racist . yall dumb
romanakudryash4|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
romanakudryash4|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
hornsby_kh|bean_colton|0.0|0.0|1.0|0.0|RT @bean_colton: Waiting in line to vote for Trump right now! #Trump2016
Amyloukingery|KamVTV|0.34|0.0|0.882|0.118|RT @KamVTV: ATTENTION TRUMP VOTERS - Here is the official Trump Voter Assistance and Ballot Security Hotline - #MyVote2016 #ElectionDay #Vo
dougsmith1946|WDFx2EU8|0.8443|0.0|0.597|0.403|"RT @WDFx2EU8:  BREAKING: WOW!!! At the last minute, Chris Matthews endorses #Trump!!! #ElectionDay  https://t.co/FjeNWIsACt"
dougsmith1946|twitter|0.8443|0.0|0.597|0.403|"RT @WDFx2EU8:  BREAKING: WOW!!! At the last minute, Chris Matthews endorses #Trump!!! #ElectionDay  https://t.co/FjeNWIsACt"
Karaszewski|twitter|0.8126|0.0|0.72|0.28|If Hillary wins we are going to drink the Blue Label... if Trump wins we are going to drink everything https://t.co/t4Sr6HnCe1
KMosetti|DRUDGE_REPORT|0.5719|0.0|0.812|0.188|@DRUDGE_REPORT @WashTimes If Mr Trump wins first thing he must do burn all of Obama executive order's.
ParkerMolloy|twitter|0.0|0.0|1.0|0.0|Team Trump mapping out the path to 270. https://t.co/C6hiikKpDW
MattJensen03|JDeezyyyy|0.0|0.0|1.0|0.0|@JDeezyyyy for trump
IMohamed2|twitter|0.0|0.0|1.0|0.0|Trump is over bud https://t.co/dVchhU2fHJ
OopsTryagain12|stevebousquet|0.4404|0.0|0.873|0.127|"RT @stevebousquet: Good news for Trump in Florida: More Republicans than Democrats are voting in Tampa Bay Tuesday, county websites say"
casxeyy|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
helovedmemore|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
helovedmemore|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
TLVRP_Tennessee|oakridger|0.1027|0.117|0.748|0.136|#Tennessee #Memphis #Nashville Trump spent a good portion of Election Day sowing doubt about the legitimacy of the https://t.co/fy868izwPk
odetosleepydun|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
odetosleepydun|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
stonesradiotx|mitchellvii|0.4404|0.0|0.838|0.162|"RT @mitchellvii: If Trump ends up dramatically outperfroming his RCP averages in early states, good sign."
X5MSport15|Pamela_Moore13|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
X5MSport15|twitter|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
1isten_up|GagePait|-0.516|0.132|0.868|0.0|RT @GagePait: #ElectionDay SHOCK EXIT POLLS:Trump up 2.3% in FlTrump up 1.2% in PaTrump up 5.3% in OhTrump up 0.8% in MichTrump up 1
xisbethprettyx|yvetteposts|0.0|0.0|1.0|0.0|RT @yvetteposts: for the 20% of the latinos voting for trump: ya moms a hoe https://t.co/SIsGBxji1L
xisbethprettyx|twitter|0.0|0.0|1.0|0.0|RT @yvetteposts: for the 20% of the latinos voting for trump: ya moms a hoe https://t.co/SIsGBxji1L
jacksonrichman|NKingofDC|-0.128|0.061|0.939|0.0|"RT @NKingofDC: So far, digging through the exits, and with the first polls about to close, there aren't a lot of signs of a looming Trump u"
LaurenDancer17|DanScavino|0.0|0.0|1.0|0.0|RT @DanScavino: Trump Campaign Headquarters-'TOP CANDIDATE QUALITY: CAN BRING CHANGE:TRUMP: 82%CLINTON: 13%#iVoted #ElectionNight #MAGA
Bscanosu21|ringer|0.0|0.0|1.0|0.0|"RT @ringer: Remember during the first debate when Trump kept telling everyone to ask Hannity, and we did? https://t.co/IEqyE0GLpH"
Bscanosu21|twitter|0.0|0.0|1.0|0.0|"RT @ringer: Remember during the first debate when Trump kept telling everyone to ask Hannity, and we did? https://t.co/IEqyE0GLpH"
rikayla|MeanwhileinCana|0.0|0.0|1.0|0.0|RT @MeanwhileinCana: #MeanwhileinCanada If Trump wins...#ElectionNight https://t.co/0dCRguut72
rikayla|twitter|0.0|0.0|1.0|0.0|RT @MeanwhileinCana: #MeanwhileinCanada If Trump wins...#ElectionNight https://t.co/0dCRguut72
mariadolderr|_thomas_27|-0.5574|0.286|0.714|0.0|@_thomas_27 not one more if you keep favoriting trump shit
ChobanianLouise|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
ChobanianLouise|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
sacapuntant|localblactivist|0.0|0.0|1.0|0.0|"RT @localblactivist: First, let's compare the obvious; Donald Trump as President Snow. https://t.co/7d62DPmIAl"
sacapuntant|twitter|0.0|0.0|1.0|0.0|"RT @localblactivist: First, let's compare the obvious; Donald Trump as President Snow. https://t.co/7d62DPmIAl"
SanpakuChi|YouTube|-0.0772|0.098|0.902|0.0|https://t.co/PXFHtx0GCx  #ElectionDay #VoteTrump - Robert De Niro exposed by Donald Trump https://t.co/N9f20yqlko via @YouTube
SanpakuChi|vote|-0.0772|0.098|0.902|0.0|https://t.co/PXFHtx0GCx  #ElectionDay #VoteTrump - Robert De Niro exposed by Donald Trump https://t.co/N9f20yqlko via @YouTube
illyahkuryahkin|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
hugva3|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
paintedtigers|DaRealDanBaulch|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
paintedtigers|t|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
hxrrera13|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Jellybean4Trump|TheDonaldNews|0.7034|0.0|0.788|0.212|RT @TheDonaldNews: LOOKING GREAT FOR @realDonaldTrump Information Showing TRUMP Up 65% in EXIT POLLS FLORIDA #FoxNews #Hannity #CNN https:/
Jellybean4Trump||0.7034|0.0|0.788|0.212|RT @TheDonaldNews: LOOKING GREAT FOR @realDonaldTrump Information Showing TRUMP Up 65% in EXIT POLLS FLORIDA #FoxNews #Hannity #CNN https:/
memeswearmatty|letters2donald|0.0|0.0|1.0|0.0|"RT @letters2donald: Children's letters to Donald Trump:  Actually, you are the snake.Violet A., age 9"
belladamaxx_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
kapustinastepa4|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
kapustinastepa4|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
zaharovfadei95|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
zaharovfadei95|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
tired_n_crabby|Thomas1774Paine|-0.3612|0.122|0.878|0.0|RT @Thomas1774Paine: #Trump Voters Complain Their Votes Locked Out of Electronic Voting Machines in New York **RT**RT**RT** #voterfraud htt
Ennio05|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: 90% of America does not approve of Congress &amp; Washington DC. Trump will DRAIN THE SWAMP! #MAGA
paulrlanni|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
m_barraza_|reIatabIe|0.0|0.0|1.0|0.0|RT @reIatabIe: Goodmorning to everyone except Donald Trump
LyndaJoHunt|jaynordlinger|0.7579|0.0|0.745|0.255|"RT @jaynordlinger: Hillary = luckiest politician ever. I know the hour is late, but are we SURE that Trump was not a Clinton plant?"
AllLivesMtr81|TallahForTrump|0.34|0.098|0.748|0.154|"RT @TallahForTrump: While KKKlinton called us Black folk Super Predators, Trump was fighting for our rights against segregation in his hote"
schul47|FrenchForTrump|0.7058|0.0|0.796|0.204|RT @FrenchForTrump: FOR THE FIRST TIME IN MY LIFEAS A FRENCH EXPATRIATEI'M SO PROUD TO CAST MY VOTEFOR DONALD J. TRUMP#ElectionDay#Vo
davidmcinnes92|Magnus_Jamieson|0.0|0.0|1.0|0.0|RT @Magnus_Jamieson: Clackmannanshire already declaring for Trump #ElectionNight
AmerPride777|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
NadineORegan|MsAmyHerron|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
NadineORegan|theguardian|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
TrumpWithUSA|JoeFreedomLove|-0.4588|0.2|0.8|0.0|RT @JoeFreedomLove: Nevada Poll Workers Break Law: Caught Wearing 'Defeat Trump' T-Shirts https://t.co/XLE9PFiyQ9
TrumpWithUSA|thegatewaypundit|-0.4588|0.2|0.8|0.0|RT @JoeFreedomLove: Nevada Poll Workers Break Law: Caught Wearing 'Defeat Trump' T-Shirts https://t.co/XLE9PFiyQ9
carradinempire|reeceking_|-0.7801|0.334|0.58|0.086|RT @reeceking_: i'm personally not focusing on putting out hella negative energy based around trump cause i don't want a negative outcome s
mks2101|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
mks2101|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
gabbie_4223|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
kdunnachie|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
fortymileFrank|fernacarieles|0.6523|0.1|0.651|0.249|"RT @fernacarieles: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://"
fortymileFrank||0.6523|0.1|0.651|0.249|"RT @fernacarieles: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://"
DSmooth_seven17|Call4AMedic|0.25|0.067|0.827|0.106|"RT @Call4AMedic: 97% of black voters are non-trump voters, again proving that black people are seriously the only smart people left among us"
linzilouxxx|AngrySalmond|-0.2944|0.153|0.744|0.103|RT @AngrySalmond: Voting for Donald Trump is a bit like deliberately infecting yourself with an STD. It's just fucking stupid. #Presidentia
RM3Barcelona4|Chappynash|-0.6705|0.234|0.766|0.0|"RT @Chappynash: @SamWiseSW Hillary is worse.  She will flip the SCOTUS into a legislative judiciary for a generation. Trump is a jerk, she"
stairwaylover|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
stairwaylover|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
greenlawley|lovelaurenxjenn|0.5719|0.0|0.821|0.179|RT @lovelaurenxjenn: If Trump or Hillary  Wins The Election I Am Moving  Out Of The Country  Goodbye America  Hello   N
thepoliticalcat|AlGiordano|0.1111|0.098|0.786|0.115|RT @AlGiordano: SPOILER ALERT: Florida votes for Clinton have already surpassed Obama 2012 as of 5 p.m. Trump lags behind Romney's. Any que
old_put|Vote3Fortrump|-0.4588|0.188|0.813|0.0|RT @Vote3Fortrump: Nevada Poll Workers Break Law: Caught Wearing Defeat Trump T-Shirts https://t.co/FKOm5pcGyI https://t.co/pAoZ6Fz2kJ
old_put|jewsnews|-0.4588|0.188|0.813|0.0|RT @Vote3Fortrump: Nevada Poll Workers Break Law: Caught Wearing Defeat Trump T-Shirts https://t.co/FKOm5pcGyI https://t.co/pAoZ6Fz2kJ
peaceharmony16|Vets_Vs_Trump|0.7404|0.0|0.77|0.23|@Vets_Vs_Trump @PAMsLOvE @MorganLsneed YOU SURE CAN BREAK THE LAW AND GET AWAY FROM IT LIKE HILLARY . THAT IS WHAT YOU ARE GOING FOR
KylanWWatson|RawStory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
KylanWWatson|rawstory|0.2732|0.0|0.851|0.149|RT @RawStory: Trump supporter pepper sprays voter at Florida polling location https://t.co/AMzlOGiAPE https://t.co/pwXo7rftEI
KaceyIlliot1669|jaketapper|-0.8687|0.376|0.542|0.081|"@jaketapper Trump is the only choice for us! Hillary cheats, lies and steals. She even cheated at the debates with help from CNN"
dronerecovery|dronerecovery|0.3182|0.0|0.859|0.141|"RT @dronerecovery: @neko_designer @ShimermanArmin ""please see the treatment of trump"" Appeal to hypocrisy, second count."
PrincessRayvXo|alyssanicholle_|0.6597|0.0|0.795|0.205|"RT @alyssanicholle_: If you vote Trump today, make sure to explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
yoAustinn|CloudN9neSyrup|0.5719|0.0|0.866|0.134|"@CloudN9neSyrup they made them for trump too, they just wait till the elections over to see who wins, and those are the ones they sell..."
NikonovFinogen|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
NikonovFinogen|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
paulaakpan|CalumSPlath|-0.6249|0.163|0.837|0.0|RT @CalumSPlath: the worst thing about a Trump presidency would be that Green Day would feel they've been given license to release another
karintracy|everywhereist|0.0|0.0|1.0|0.0|"@everywhereist @jasonvolack @ABC If I were #Trump, I would stuff the baker here. Ye gads..."
mi4of5jaa|BruceBartlett|0.6311|0.076|0.688|0.235|"RT @BruceBartlett: For the record, I voted enthusiastically for Hillary Clinton today. She may not be perfect, but she's light years better"
andreablu_it|goldengateblond|-0.7184|0.222|0.778|0.0|RT @goldengateblond: The Trump campaign asked a judge to make the names of Nevada poll workers public. She had no time for their bullshit.
Mrgee_bande|Ary_AntiPT|0.0|0.0|1.0|0.0|"RT @Ary_AntiPT: Trump up 70.5% to Hillary's 25.8% in Indiana. 35,646 votes to 13,049 #ElectionNight"
charliewalton11|YouTube|0.5267|0.0|0.746|0.254|Final Electoral College Map Trump is winning November 8 https://t.co/h9Ie0Mjgcq via @YouTube
charliewalton11|youtube|0.5267|0.0|0.746|0.254|Final Electoral College Map Trump is winning November 8 https://t.co/h9Ie0Mjgcq via @YouTube
1965Randy|youtube|0.0|0.0|1.0|0.0|Donald trumps song for his hair  https://t.co/yYa1VRuGgH  #ElectionNight #Trump #Trump2016  #trump
timofeevbonifa3|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
timofeevbonifa3|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
RenaldIgnatov|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
RenaldIgnatov|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
esmerugh|CherOfficiaI|0.6633|0.0|0.783|0.217|RT @CherOfficiaI: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
tommyshida|staffsgtshawnb2|0.5267|0.0|0.726|0.274|RT @staffsgtshawnb2: #FoxNews2016.  trump is winning new Hampshire. 52 41
jonathancristol|jaynordlinger|0.4404|0.0|0.884|0.116|RT @jaynordlinger: If Bill Clinton talked Donald Trump into running for the GOP nomination -- Clinton truly is the wiliest politician in wo
NathanTunell|goldengateblond|-0.7184|0.222|0.778|0.0|RT @goldengateblond: The Trump campaign asked a judge to make the names of Nevada poll workers public. She had no time for their bullshit.
Donnalee711|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
TsayPA|chrislhayes|0.0|0.0|1.0|0.0|"RT @chrislhayes: After waiting until almost *literally* the last moment, Toomey votes and says he voted for Trump."
Gingerbreadhau5|Thomas_A_Moore|0.0|0.0|1.0|0.0|RT @Thomas_A_Moore: how it feels to vote against Trump https://t.co/9oy8jsjtv3
Gingerbreadhau5|twitter|0.0|0.0|1.0|0.0|RT @Thomas_A_Moore: how it feels to vote against Trump https://t.co/9oy8jsjtv3
diva6684|MSignorile|-0.8481|0.349|0.586|0.065|RT @MSignorile: Trump &amp; GOP are putting gun to Americas head: Elect #Trump or we create complete havoc. Dont fall for threats. Stop them.
Cato_Cat|peddoc63|0.3182|0.0|0.905|0.095|"RT @peddoc63: My 19 year old son 1st supported Bernie Sanders, then Gary Johnson, today he is voting for Donald J. Trump#ElectionNight #m"
XicanoAdrian|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
XicanoAdrian|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
niallsayspotato|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
niallsayspotato|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
theOGericmullin|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
neanybean18|sweetatertot2|0.0|0.0|1.0|0.0|RT @sweetatertot2: Florida residents we need you head to the polls &amp; #Vote2016 for Trump. Florida is needed! #ElectionDay #Election2016 #WT
sobercat13|FoxBusiness|0.8283|0.201|0.429|0.37|@FoxBusiness PLEASE STOP WHINING. The numbers are not in &amp; you are all ready finding people to blame. Trump got GREAT FREE network coverage!
SetarehSabety|facebook|0.0|0.0|1.0|0.0|Here we go... Trump candidacy collateral damage... #electionday Where the h is Azusa? https://t.co/2jdzUsMd3O
DawnShmawn|AnnCoulter|-0.5106|0.13|0.87|0.0|"@AnnCoulter  meanwhile since the rise of Donald trump the KKK is handing out fliers again and hanging black people. Ann, you're an idiot."
lkinglwt|justinalvarez98|0.691|0.0|0.725|0.275|RT @justinalvarez98: Honestly if you voted for Trump unfollow me I don't need that negativity in my life.
burova_aleksa|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
burova_aleksa|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
bjstatha|0hour|0.0|0.0|1.0|0.0|RT @0hour: Everyone grab your Cell phones call people and get more votes!TRUMPGO GO GO! https://t.co/tNqo6MPUT5
bjstatha|twitter|0.0|0.0|1.0|0.0|RT @0hour: Everyone grab your Cell phones call people and get more votes!TRUMPGO GO GO! https://t.co/tNqo6MPUT5
She_is_morg|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
She_is_morg|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
dailycosmic|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: 90% of America does not approve of Congress &amp; Washington DC. Trump will DRAIN THE SWAMP! #MAGA
Battleborne|realDonaldTrump|0.6037|0.0|0.696|0.304|#FoxNews2016.@realDonaldTrump  #Election2016 Results: NH 1% rpt Trump 52% Clinton 41%
Andulos|conservativluke|0.0|0.0|1.0|0.0|@conservativluke @waynedupreeshow Ah my apologies then. I guess I'm just too used to seeing Trump's hitler youth.
EceeR___|ImageSlays|-0.1531|0.096|0.904|0.0|RT @ImageSlays: If Donald Trump Looses the election I'll give everybody who RTs this $5 PayPal.
caaroliinam|OliviaMesser|0.6124|0.0|0.5|0.5|"RT @OliviaMesser: Like father, like son:https://t.co/HjNUN2POX9 https://t.co/ToamX6hNk0"
caaroliinam|thedailybeast|0.6124|0.0|0.5|0.5|"RT @OliviaMesser: Like father, like son:https://t.co/HjNUN2POX9 https://t.co/ToamX6hNk0"
DattNigga_Quan|DaRealGleesh|-0.5423|0.467|0.533|0.0|RT @DaRealGleesh: Fuck Donald trump 
ChpaMaud|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
ChpaMaud|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
lmanzanillad|PpollingNumbers|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
lmanzanillad|twitter|0.0|0.0|1.0|0.0|RT @PpollingNumbers: Final @trfgrp Electoral Map(270 EV Needed):Trump 306Clinton 232 https://t.co/Kf3IaODMhD
Pas_Normal|TBNSport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
Pas_Normal|tbnsport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
C_Wade21|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
C_Wade21|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
BatflecksRobin|EmilyBett|0.4404|0.0|0.508|0.492|@EmilyBett trump is better
Heckel_n_Jeckel|0hour|0.0|0.0|1.0|0.0|RT @0hour: Paris Hilton voted Trump BTFO!
OfNannaAndMen|jaw_cee|0.431|0.0|0.898|0.102|RT @jaw_cee: If you're Mexican &amp; voting for Trump let me just say: 1. He doesn't give a fuck about you2. Eres un pendejo3. We don't clai
JimbauxsJournal|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
JimbauxsJournal|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
ScottTh24545752|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
ScottTh24545752|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
maritundra|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
maritundra|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
Jennife51072808|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
snugglebutt21|dril|-0.7845|0.264|0.736|0.0|RT @dril: donlad trump reportedly says that normal type pokemon are a waste of time. they're just dirty birds &amp; rats who have no right bein
BballShizzle|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
BballShizzle|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
bigstewo7|yankeebrit77|0.4215|0.0|0.887|0.113|"@yankeebrit77 @Pamela_Moore13 nice how they say "" they try to vote for one candidate, just to have their vote switch to another"" only trump"
ggullotti1|Miikeyyv|-0.3476|0.186|0.814|0.0|@Miikeyyv @DlCKFORD @jojo_bear32 @jackwilsonnnnnn liberals don't understand the value of hard work. They depend on handouts #Trump
Mapada1|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
Mapada1|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
Kike_Loves_LA14|YG|-0.5719|0.371|0.479|0.15|"RT @YG: All trump supports unfollow me, &amp; Suck my dick"
E46lopez|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
E46lopez|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
paniela100|alaskantexanQCT|0.0|0.0|1.0|0.0|RT @alaskantexanQCT: Yo fam heading to Philly with some homies and 2 vans. Gonna take Black Trump voters 2 the polls ALL DAY tomorrow! #MAG
ljwnorth|BBCWillVernon|0.4019|0.0|0.828|0.172|"RT @BBCWillVernon: Pro-Trump Russian politicians, activists, journalists at a US #ElectionNight party in #Moscow https://t.co/iV2UN65aFY"
ljwnorth|twitter|0.4019|0.0|0.828|0.172|"RT @BBCWillVernon: Pro-Trump Russian politicians, activists, journalists at a US #ElectionNight party in #Moscow https://t.co/iV2UN65aFY"
TLVRP_Tennessee|wmcactionnews5|0.0|0.0|1.0|0.0|"#Tennessee #Memphis #Nashville Finally, it's Clinton or Trump: Long race ends, voters pick https://t.co/8rt7Kr4Upu"
creminsmom|MCrisCardena|-0.4003|0.119|0.881|0.0|@MCrisCardena If Hillary worked for a bank (any US Company) &amp;  released Confidential Info.... She is fired.... Fire Hillary .... Vote Trump!
NormandinRob|trump_florida|0.4019|0.0|0.828|0.172|RT @trump_florida: Source: The Military Times951 Active Duty Troops PolledTrump 54%     Hillary 25%#TrumpPence16 https://t.co/t1n374qx7M
NormandinRob|twitter|0.4019|0.0|0.828|0.172|RT @trump_florida: Source: The Military Times951 Active Duty Troops PolledTrump 54%     Hillary 25%#TrumpPence16 https://t.co/t1n374qx7M
biebertopping|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
biebertopping|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
Republican1950|jerome_corsi|0.1591|0.066|0.844|0.089|RT @jerome_corsi: Lines in many states are LONG - BE RESOLVED TO STAY IN LINE until you get to VOTE FOR TRUMP - nothing is more important t
TrailKing71|kayleighmcenany|0.7177|0.0|0.769|0.231|"RT @kayleighmcenany: Trump has a .2% lead in Florida according to Real Clear Politics. My fellow Floridians, get out, vote, &amp; take friends!"
rmcardz|0hour|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
rmcardz|twitter|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
noukanat|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
kelsheintz|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
kelsheintz|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
_Dobbins_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
PaulMakesMovies|TIME|0.4019|0.0|0.856|0.144|RT @TIME: Mixed Drinks are $13 and beer is $11 at Donald Trump's election night party https://t.co/GqEEQDeBCf
PaulMakesMovies|fortune|0.4019|0.0|0.856|0.144|RT @TIME: Mixed Drinks are $13 and beer is $11 at Donald Trump's election night party https://t.co/GqEEQDeBCf
samsgotskills|Cain_Unable|0.0|0.0|1.0|0.0|"RT @Cain_Unable: I just tried to Vote Trump &amp; the staff wouldn't let me just because I'm ""in Kent"" &amp; ""this is a Tesco self service checkout"
emastiffs|PeterSweden7|0.0|0.0|1.0|0.0|"RT @PeterSweden7: So far with votes counted in IN, KY &amp; NH:Trump: 149 808 (68%)Clinton: 62 250 (28%)#ElectionNight"
Healyjauregay|fifthorgajsms|0.0|0.0|1.0|0.0|RT @fifthorgajsms: Mexicans/gays/latinos/blacks/women for Trump!!! Me:#ElectionDay https://t.co/OKlNr5Da5u
Healyjauregay|twitter|0.0|0.0|1.0|0.0|RT @fifthorgajsms: Mexicans/gays/latinos/blacks/women for Trump!!! Me:#ElectionDay https://t.co/OKlNr5Da5u
cbest00|twitter|0.0|0.0|1.0|0.0|TRUMP https://t.co/EdduLFrePc
haleylujaaah|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
CocoRoberts2|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: Right now, Trump is making up more than half of Obama's entire 2012 margin of victory in FL in JUST ONE COUNTY!"
Mr_NastyTime623|castle2410|-0.763|0.376|0.501|0.123|@castle2410 We really really hate him down here.....more than Trump...now he's definitely a known racist
feeIingmyoats|melaninbarbie|-0.8481|0.286|0.714|0.0|"RT @melaninbarbie: Any black person that votes for Trump gets last pick for shade spots. If you get a dead bush with no leaves, too damn ba"
Ontapron|mitchellvii|0.2177|0.137|0.684|0.179|RT @mitchellvii: So was Trump winning CO and conveniently every voting machine in the state broke?
hwomack2525|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
birdlady19492|mitchellvii|0.7998|0.0|0.736|0.264|RT @mitchellvii: The last RCP Poll had Trump winning KY by 17.  He is currently winning by 52 points.Monster vote?  Dem crossovers?
rldods|realDonaldTrump!|0.0|0.0|1.0|0.0|I am going to go ahead call #Georgia for @realDonaldTrump! #Trump earns 16 #electoralvotes @WorthItElection
Jleitner7|TheFunnyVine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
Jleitner7|vine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
PileOfSierra|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
PileOfSierra|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
rabuliz|DonaldJTrumpJr|0.9059|0.0|0.394|0.606|RT @DonaldJTrumpJr: Thank you! Love the energy and enthusiasm! #MAGA #Trump https://t.co/MZfYawGs5l
rabuliz|twitter|0.9059|0.0|0.394|0.606|RT @DonaldJTrumpJr: Thank you! Love the energy and enthusiasm! #MAGA #Trump https://t.co/MZfYawGs5l
jackalate|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
buttonlol|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
alison8796|Variety|0.0|0.0|1.0|0.0|RT @Variety: George W. Bush didn't vote for Donald Trump or Hillary Clinton for president https://t.co/JaXKzBWOTY https://t.co/CspXjAF5AS
alison8796|variety|0.0|0.0|1.0|0.0|RT @Variety: George W. Bush didn't vote for Donald Trump or Hillary Clinton for president https://t.co/JaXKzBWOTY https://t.co/CspXjAF5AS
ponomarevaippo6|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ponomarevaippo6|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
CHOCLABLOVER|azmoderate|-0.5267|0.313|0.568|0.119|RT @azmoderate: Trump supporter arrested after pulling gun at Florida polling station https://t.co/uK8MC3TKqX
CHOCLABLOVER|rawstory|-0.5267|0.313|0.568|0.119|RT @azmoderate: Trump supporter arrested after pulling gun at Florida polling station https://t.co/uK8MC3TKqX
The_Walz|twitter|0.6249|0.0|0.702|0.298|"Prediction 1: Trump does well, but not enough. This is the safest bet. https://t.co/8stIga1eLC"
MatJoseph1|DonaldJTrumpJr|0.6739|0.0|0.688|0.312|@DonaldJTrumpJr @realDonaldTrump PRESIDENT DONALD J TRUMP WILL BE THE WINNER TONIGHT. #MAKEHILARYCLINTONCRY
GoinsteadySki|JohnJohnDaDon|0.0|0.0|1.0|0.0|RT @JohnJohnDaDon: Just cuz you Anti-Trump doesn't mean you have to be Pro-ClintonEspecially if you're considered a minority
Tvirden09|PolitixGal|0.1779|0.101|0.769|0.13|"RT @PolitixGal: TRUMP --&gt; The man that gave up his billionaire lifestyle to be ridiculed, slandered &amp; mistreated to save America."
schmemmm|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
schmemmm|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
kulikovbesson|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
kulikovbesson|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
Only_Oneydi|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
kentran65|michellerj1019|0.0|0.0|1.0|0.0|"RT @michellerj1019: Trump leads Clinton by 120,000 votes  the first Republican candidate to EVER lead in early voting in Florida. #Electio"
Cinemadreams_|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
Cinemadreams_|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
diodoraaksyono3|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
diodoraaksyono3|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
Princesstoe|ENuFFZnuFF2001|0.5904|0.0|0.723|0.277|RT @ENuFFZnuFF2001: TRUMP NEEDS FLORIDA CALL YOUR FRIENDS VOTE VOTE https://t.co/jeK3ro5Gqw
Princesstoe|twitter|0.5904|0.0|0.723|0.277|RT @ENuFFZnuFF2001: TRUMP NEEDS FLORIDA CALL YOUR FRIENDS VOTE VOTE https://t.co/jeK3ro5Gqw
korbyn00|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
TimGclaw|sturdyAlex|-0.228|0.091|0.909|0.0|RT @sturdyAlex: The Trump men appear a little worried about the female vote. Including that of their wives. (h/t @durrant_james) https://t.
TimGclaw||-0.228|0.091|0.909|0.0|RT @sturdyAlex: The Trump men appear a little worried about the female vote. Including that of their wives. (h/t @durrant_james) https://t.
MoneyMills_72|garrettrt21|0.1901|0.0|0.889|0.111|RT @garrettrt21: I like how my snapchat has the trump filter but not the Hilary one#TrumpTrain
Gibbe84|rblandford|-0.5574|0.31|0.69|0.0|RT @rblandford: Shit. Sunderland South have gone for Trump.
terrydvl|theglobaluniter|0.0|0.0|1.0|0.0|RT @theglobaluniter: If you live in the Panhandle area of Florida we need you to go and #Vote #Trump.A call to action by .@DonaldJTrumpJ
DevloPM|SoaRPraizist|0.5719|0.0|0.802|0.198|"RT @SoaRPraizist: If Trump wins the election, I will make artwork for everyone that RTs this tweet"
dancodesigns|jasonvolack|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
dancodesigns|twitter|0.0|0.0|1.0|0.0|RT @jasonvolack: A Donald Trump cake being wheeled into Trump Tower @abc #ElectionDay https://t.co/HSkHChfUSA
TheKStainback|pattymo|0.0772|0.0|0.936|0.064|"RT @pattymo: BAKER: Hey, what kind of expression do you want on his faceTRUMP STAFFER: Let's go with ""haunted"" https://t.co/SxNJQX4r2F"
TheKStainback|twitter|0.0772|0.0|0.936|0.064|"RT @pattymo: BAKER: Hey, what kind of expression do you want on his faceTRUMP STAFFER: Let's go with ""haunted"" https://t.co/SxNJQX4r2F"
allanktbh|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
shouldbenow|Houseman75|0.5574|0.0|0.806|0.194|RT @Houseman75: I proudly and unequivocally voted for Donald J. Trump for President. #FoxNews2016 #TrumpPence16 #SaveTheCoalMiner https://t
shouldbenow||0.5574|0.0|0.806|0.194|RT @Houseman75: I proudly and unequivocally voted for Donald J. Trump for President. #FoxNews2016 #TrumpPence16 #SaveTheCoalMiner https://t
RaulAriasZamor2|AmericasVoice|-0.2023|0.094|0.848|0.058|RT @AmericasVoice: BREAKING: National exit poll number for Latino Voters from @LatinoDecisions: Clinton 79 - Trump 18. New low for GOP. Sam
teakinrj|thinkprogress|0.0|0.0|1.0|0.0|RT @thinkprogress: Drawing out voters of color in Trump territory https://t.co/WR6kFMtK17 #ElectionDay https://t.co/rkFoUbECHj
teakinrj|medium|0.0|0.0|1.0|0.0|RT @thinkprogress: Drawing out voters of color in Trump territory https://t.co/WR6kFMtK17 #ElectionDay https://t.co/rkFoUbECHj
SAILORSOLEMN|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
TracyB80484834|HillaryClinton|0.128|0.177|0.622|0.201|"RT @HillaryClinton: Today, let's show the world that love will always trump hate. https://t.co/jfd3CXu1CS https://t.co/a7FXGtAfiG"
TracyB80484834|hillaryclinton|0.128|0.177|0.622|0.201|"RT @HillaryClinton: Today, let's show the world that love will always trump hate. https://t.co/jfd3CXu1CS https://t.co/a7FXGtAfiG"
dcwishy|JOMainEvent|0.7081|0.0|0.754|0.246|"RT @JOMainEvent: I don't know about you guys, but this is crucial! We all know Trump supporters want Change!#ElectionNight #voted #TeamT"
SomeGuysCat|alcardfan|0.296|0.0|0.896|0.104|RT @alcardfan: I voted for Donald Trump and Mike Pence. Will you join me? Find your polling place: https://t.co/N8aoPrumfM #TrumpTrain #Ele
SomeGuysCat|vote|0.296|0.0|0.896|0.104|RT @alcardfan: I voted for Donald Trump and Mike Pence. Will you join me? Find your polling place: https://t.co/N8aoPrumfM #TrumpTrain #Ele
harvestlimited|DaveSilberman|0.5859|0.12|0.598|0.282|"RT @DaveSilberman: Broke out the good wine. Because, if Trump wins, what exactly am I saving it for?"
xXx_MattMan_xXx|mitchellvii|0.4648|0.0|0.664|0.336|"RT @mitchellvii: Again, HUGE FOR TRUMP. https://t.co/osXpZyBcze"
xXx_MattMan_xXx|twitter|0.4648|0.0|0.664|0.336|"RT @mitchellvii: Again, HUGE FOR TRUMP. https://t.co/osXpZyBcze"
milen_ershov|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
milen_ershov|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
vintage57|GaryLineker|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
vintage57|twitter|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
KarenTr58210895|Ocean_State211|0.0|0.0|1.0|0.0|RT @Ocean_State211: BREAKING: The first Florida exit poll numbers have been released.Trump 55%Clinton 39%Johnson 6% THIS IS A #HOAX!!
kdotkitty|JamilahLemieux|-0.2732|0.087|0.87|0.043|"RT @JamilahLemieux: No matter what happens tonight, the fact that Donald Trump has gotten this far is a stain on America that can't be wash"
JR777771|MarkJGrimaldi|0.0|0.0|1.0|0.0|RT @MarkJGrimaldi: It's official! #DonaldTrump has made history! https://t.co/j3zs41QwJ6.#TaxReturns #ImWithHer #NeverTrump #ElectionDay #
JR777771|t|0.0|0.0|1.0|0.0|RT @MarkJGrimaldi: It's official! #DonaldTrump has made history! https://t.co/j3zs41QwJ6.#TaxReturns #ImWithHer #NeverTrump #ElectionDay #
basedruba|dj_rocklee|0.5374|0.082|0.752|0.166|RT @dj_rocklee: Shiiitttt if Donald Trump wins this election im warning ALL YALL !!!!! Knuck if you buck white America. Knuck if you the
Colville|Daniel_Ohana|0.7177|0.0|0.6|0.4|RT @Daniel_Ohana: Electrify your Trump sign for instant justice! :-) https://t.co/jHSUqbFz0Q
Colville|twitter|0.7177|0.0|0.6|0.4|RT @Daniel_Ohana: Electrify your Trump sign for instant justice! :-) https://t.co/jHSUqbFz0Q
UnicornsSA|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
coconutbih|1942bs|0.6339|0.082|0.65|0.268|RT @1942bs: don't you dare disrespect Michael Jackson like this. He would not support a Trump as a politician if he were alive https://t.co
coconutbih|t|0.6339|0.082|0.65|0.268|RT @1942bs: don't you dare disrespect Michael Jackson like this. He would not support a Trump as a politician if he were alive https://t.co
bethjan5|realDonaldTrump|0.68|0.0|0.752|0.248|"@realDonaldTrump Thank you Mr. Trump, you've done more for America than you know.  All our hopes are with you!"
avenira_yudina|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
avenira_yudina|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
graememurphy77|HalleyBorderCol|0.0|0.0|1.0|0.0|RT @HalleyBorderCol: KY @ 4% reporting hasTrump 66Crooked 29THIS IS BIGPolls had Trump at +17#MAGA!
SandieHelm|BarbMuenchen|0.4796|0.0|0.865|0.135|RT @BarbMuenchen: URGENT! Calling all #Florida voters and PanHandle of #Florida voters Get out and vote! Trump campaign calling all voters
WoodJustRuff|FantasyDouche|-0.6486|0.212|0.788|0.0|"RT @FantasyDouche: If Donald Jr. and Eric Trump go to Westworld, what's the over/under on dead hookers?"
SaraWillingham2|Jace51Jm|0.0|0.0|1.0|0.0|RT @Jace51Jm: King Trump! https://t.co/vrQ6GQWBS2
SaraWillingham2|twitter|0.0|0.0|1.0|0.0|RT @Jace51Jm: King Trump! https://t.co/vrQ6GQWBS2
JoshNoneYaBiz|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
JoshNoneYaBiz|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
summeeriynn|HoodBibIe|0.3612|0.082|0.781|0.138|RT @HoodBibIe: Stop saying if trump wins yall moving out of the country.  Stfu yall cant even move outta ya mommas house https://t.co/k
summeeriynn|twitter|0.3612|0.082|0.781|0.138|RT @HoodBibIe: Stop saying if trump wins yall moving out of the country.  Stfu yall cant even move outta ya mommas house https://t.co/k
friwaysblog|costareports|0.0|0.0|1.0|0.0|"RT @costareports: On the phone w/ Giuliani. He just left Trump's apt. Said Trump is ""watching everything even tho I'm telling him not to."""
CLEFAlRlES|drewtoothpaste|0.4215|0.0|0.865|0.135|RT @drewtoothpaste: ME: anyone but trumpGARY JOHNSON: I will outlaw schools.JILL STEIN: Crystals are the only technology we need.ME: ok
fordstokes|KarlRove|-0.4767|0.307|0.693|0.0|@KarlRove Unfair shot at Trump on Election night.
lainied_|brooke_hawley5|0.0|0.0|1.0|0.0|RT @brooke_hawley5: Cant wait until Barack Obama is finally out of office tomorrow and Donald Trump is our next precedent #MakeAmericaGrea
ThomasAHester2|spkhp|-0.0516|0.134|0.741|0.125|"RT @spkhp: Me: what do you know about Donald trumpKinder: Donald Trump hates Black peopleMe: Hmm, interesting https://t.co/8dMLIuUWg4"
ThomasAHester2|twitter|-0.0516|0.134|0.741|0.125|"RT @spkhp: Me: what do you know about Donald trumpKinder: Donald Trump hates Black peopleMe: Hmm, interesting https://t.co/8dMLIuUWg4"
JohnnyMooor|FunnyPicsDepot|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
JohnnyMooor|twitter|0.8126|0.0|0.575|0.425|RT @FunnyPicsDepot: Me if Trump wins vs. Me if Hilary wins https://t.co/Ghqdn4X7Cv
SaintCarolyn6|dmckinney218|0.0|0.0|1.0|0.0|RT @dmckinney218: Pennsylvania voting for Donald Trump! https://t.co/4iRP2RH0Jz
SaintCarolyn6|twitter|0.0|0.0|1.0|0.0|RT @dmckinney218: Pennsylvania voting for Donald Trump! https://t.co/4iRP2RH0Jz
JenniferDonels2|LVonrobke|0.8777|0.0|0.675|0.325|RT @LVonrobke: We voted to make America great again ! #TrumpPence16  Thank you Mr Trump for all you do and for caring about middle America
gordon1470|realDonaldTrump|0.9285|0.0|0.542|0.458|RT @realDonaldTrump: Happy #CincoDeMayo! The best taco bowls are made in Trump Tower Grill. I love Hispanics! https://t.co/ufoTeQd8yA https
gordon1470|facebook|0.9285|0.0|0.542|0.458|RT @realDonaldTrump: Happy #CincoDeMayo! The best taco bowls are made in Trump Tower Grill. I love Hispanics! https://t.co/ufoTeQd8yA https
steve62269|cristinalaila1|0.0|0.0|1.0|0.0|RT @cristinalaila1: Just waited 45 minutes in line and voted for Trump #MAGA3X #MAGASelfie #ElectionDay2016 #MyVote2016 https://t.co/c0
steve62269|t|0.0|0.0|1.0|0.0|RT @cristinalaila1: Just waited 45 minutes in line and voted for Trump #MAGA3X #MAGASelfie #ElectionDay2016 #MyVote2016 https://t.co/c0
payge_14|Peifer21|0.0|0.0|1.0|0.0|RT @Peifer21: All of you sheep minded idiots/frauds can go f**k yourselves.  Go Trump! https://t.co/jPtPAZi9sA
payge_14|twitter|0.0|0.0|1.0|0.0|RT @Peifer21: All of you sheep minded idiots/frauds can go f**k yourselves.  Go Trump! https://t.co/jPtPAZi9sA
sitocyrus|JackJ|0.5719|0.0|0.764|0.236|@JackJ if donald trump wins i let you live in my home in spain 
aspen1031|blvckpapii|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
aspen1031|twitter|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
c_hallll|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
JulionficMy|ViraI|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
JulionficMy|twitter|-0.5213|0.187|0.813|0.0|RT @ViraI: Some voting machines will not allow you to vote for Donald Trump. They are looking into the problem. https://t.co/bh58Q7kIvT
magicbravosolo|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
elmorephd|NRO|0.0|0.0|1.0|0.0|"RT @NRO: Early Exit Polls: Trump Opens YUGE Gap between College-Educated, Non-College-Educated Whiteshttps://t.co/ADpCNhYfiC #ElectionNight"
dale_bernadette|seanhannity|-0.4574|0.187|0.813|0.0|@seanhannity Pennsylvania voters complained of their vote 2 Trump wld switch to Hillary. Frauding again?!
jackramseyy|cujoknows|0.0|0.0|1.0|0.0|RT @cujoknows: Donald Trump's electoral map taking form.... #L https://t.co/WSQeNqrQkt
jackramseyy|twitter|0.0|0.0|1.0|0.0|RT @cujoknows: Donald Trump's electoral map taking form.... #L https://t.co/WSQeNqrQkt
xora613|tpalmore|0.686|0.0|0.739|0.261|RT @tpalmore: From a military veteran!! Please go out and vote for Trump! Don't be fooled by the media!
hannnahvogel|Selmani__|0.0|0.0|1.0|0.0|RT @Selmani__: If you voted for trump your moms a hoe
Waybino|WorIdStarComedy|0.8126|0.0|0.575|0.425|RT @WorIdStarComedy: Me if Trump wins vs. Me if Hilary wins https://t.co/C7ydgHXWyQ
Waybino|twitter|0.8126|0.0|0.575|0.425|RT @WorIdStarComedy: Me if Trump wins vs. Me if Hilary wins https://t.co/C7ydgHXWyQ
seanwlknsn|aduanebrown|0.0|0.0|1.0|0.0|"RT @aduanebrown: One thing we can see: Even though it's early, Trump is over-performing his polling averages in the 2 states we have raw nu"
cjmcginnis|travelskills|0.0|0.0|1.0|0.0|"One night at the Trump International Hotel in Washington,DC https://t.co/m4NzI16Irv https://t.co/CjL9COI506"
therightworks|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
CathyLanier3|DonaldJTrumpJr|0.6705|0.0|0.792|0.208|RT @DonaldJTrumpJr: In 2000 New Mexico was determined by less than 400 votes. Every single vote counts. Your vote counts. Call your friends
Doryphonehome|CrisCovaDiaz|0.0|0.0|1.0|0.0|RT @CrisCovaDiaz: I'm also a #CollegeEducatedLatina voting specifically against Trump. @ananavarro #ElectionNight #myvote2016 https://t.co/
Doryphonehome|t|0.0|0.0|1.0|0.0|RT @CrisCovaDiaz: I'm also a #CollegeEducatedLatina voting specifically against Trump. @ananavarro #ElectionNight #myvote2016 https://t.co/
vatiammatri|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
MWatsPatriot|nbcconnecticut|0.0|0.0|1.0|0.0|#trumpI just told #NBCCT I voted today for Donald #Trump. Follow @nbcconnecticut for the latest election news. https://t.co/IX8mb1stcJ
MWatsPatriot|nbcconnecticut|0.0|0.0|1.0|0.0|#trumpI just told #NBCCT I voted today for Donald #Trump. Follow @nbcconnecticut for the latest election news. https://t.co/IX8mb1stcJ
djlithium|DonaldJTrumpJr|0.5696|0.0|0.872|0.128|"RT @DonaldJTrumpJr: If you have friends in MI, OH, FL, PA -- CALL THEM and tell them to VOTE TRUMP! You can make a difference! #MAGA #Tru"
Ripchord12|RichardGrenell|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
Ripchord12|twitter|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
tadiadunton|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
tadiadunton|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
comment_here|mitchellvii|0.7998|0.0|0.736|0.264|RT @mitchellvii: The last RCP Poll had Trump winning KY by 17.  He is currently winning by 52 points.Monster vote?  Dem crossovers?
douniahamad_|FunctionUp|0.8672|0.071|0.578|0.351|"RT @FunctionUp: Or maybe it's because Trump is a disgusting man who spews nothing but hate. But sure, teenagers hate him ""because Twitter h"
happkat|0hour|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
happkat|twitter|-0.7317|0.359|0.641|0.0|RT @0hour: REPEAT AFTER ME DONALD J TRUMP WILL BE PRESIDENT NO DOUBTS! https://t.co/FFc5B4oQE2
DeniseSWells63|JaimeeLiegh|0.8885|0.0|0.61|0.39|RT @JaimeeLiegh: pretty sure if Trump wins Europe is going to suddenly increase in population because of the amount of Americans migrating
neatIester|StanceFrac|0.5719|0.0|0.791|0.209|RT @StanceFrac: If Donald trump wins the election I'll PayPal everyone that rted this $1
Mariaebrothert2|DonaldJTrumpJr|0.6705|0.0|0.792|0.208|RT @DonaldJTrumpJr: In 2000 New Mexico was determined by less than 400 votes. Every single vote counts. Your vote counts. Call your friends
bdarlingwhite|MMFlint|0.0|0.0|1.0|0.0|RT @MMFlint: Michigan! They say it's going to be close! GO VOTE NOW! Our state has been on the ropes for years. Trump will finish us off. G
JayJay2016Mma|bakedalaska|0.4225|0.16|0.621|0.219|RT @bakedalaska: I am so proud to have voted for Donald J. Trump today. Couldn't be happier. Thank you everyone for your support. #MAGASe
tmcmill81|costareports|0.0|0.0|1.0|0.0|"RT @costareports: On the phone w/ Giuliani. He just left Trump's apt. Said Trump is ""watching everything even tho I'm telling him not to."""
iamblissss|drvixfutures|0.1027|0.165|0.692|0.142|"@drvixfutures 13s or lower, unless Trump wins. Do you remember how low UVXY went before the last reverse split? Around 6 I believe."
EwanHawking|mitchellvii|0.5719|0.0|0.85|0.15|"RT @mitchellvii: Romney won Brevard County by 36,000 votes in 2012.  I calculate Trump leads it by 52,000 votes.  +16,000 votes for Trump o"
DianaLTaub|MIGOP|-0.5411|0.253|0.658|0.089|"@MIGOP @MichiganDems @UMichFootball @realDonaldTrump okay Trumpsters , no worry dems, your allowed to vote for Trump..vote Trump now!"
dihelfrich|tinkrbel5|-0.5106|0.125|0.875|0.0|RT @tinkrbel5: @DonaldJTrumpJr @Frankhe1 Right now I am sick of the soros owned machines recording Trump votes as Hillary in PA FL CA NC &amp;
_nguwop|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
_nguwop|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
techdeckturtle|popss0n|0.0|0.0|1.0|0.0|RT @popss0n: Trump for president 
gurr_john|abkbundy|0.0|0.0|1.0|0.0|"RT @abkbundy: Trump becomes the first to break 100,000 votes tonight. #ElectionNight"
drafthorse2012|mitchellvii|0.2177|0.137|0.684|0.179|RT @mitchellvii: So was Trump winning CO and conveniently every voting machine in the state broke?
DJ_Homewrecker|DJ_Homewrecker|-0.5319|0.209|0.791|0.0|RT @DJ_Homewrecker: TRUMP IS ABOUT TO LOSE AN ELECTION ON TACO TUESDAY. SO FITTING.
MillenniumMayor|Veteran4Trump|0.4926|0.0|0.856|0.144|@Veteran4Trump @realDonaldTrump as a. Veteran my wife and I voted for Trump/Pence even though we live in California it felt good !
jabs611|TeresaEdelglass|0.471|0.0|0.839|0.161|RT @TeresaEdelglass: Voting machine in #PA refuses to allow vote for @realDonaldTrumpWe are the watchdogs!REPORT! REPORT! REPORT! h
VanessaLuver_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
VanessaLuver_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
KoolaidUSA|NewYorker|0.4588|0.0|0.842|0.158|RT @NewYorker: The Trump campaign was laughed out of the courtroom in Nevada today. https://t.co/XpavP0b3k8 #ElectionDay https://t.co/hmjmK
KoolaidUSA|newyorker|0.4588|0.0|0.842|0.158|RT @NewYorker: The Trump campaign was laughed out of the courtroom in Nevada today. https://t.co/XpavP0b3k8 #ElectionDay https://t.co/hmjmK
lonerismism|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
realSpottswoode|mitchellvii|0.7284|0.0|0.61|0.39|RT @mitchellvii: TRUMP IS GOING TO WIN!  GO VOTE!
Sayitaintdaun|twitter|0.0|0.0|1.0|0.0|Is Hillary and Trump running still? https://t.co/13E4XJNOvo
tayb7|Storyteller1951|0.0|0.0|1.0|0.0|"RT @Storyteller1951: ""@KYWrangler: Voted in KY! #MAGASELFIE @MAGA3X @Cernovich @realDonaldTrump https://t.co/BGXzbM6M6Q"" Vote Trump watch o"
tayb7|twitter|0.0|0.0|1.0|0.0|"RT @Storyteller1951: ""@KYWrangler: Voted in KY! #MAGASELFIE @MAGA3X @Cernovich @realDonaldTrump https://t.co/BGXzbM6M6Q"" Vote Trump watch o"
ranpaq|HalleyBorderCol|0.7703|0.0|0.74|0.26|"RT @HalleyBorderCol: For anyone wanting election results as them come in, the Guardian site seems quite good. Looking good for #Trump!htt"
pmswolfy|cook_jengle|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
pmswolfy|twitter|0.0|0.0|1.0|0.0|RT @cook_jengle: #Election2016 Voted for Trump! https://t.co/n2YXWve3qm
GelasiyKuzmin|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
GelasiyKuzmin|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ilhaanxo|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
Lurvsammx|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
nschim|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
koalagirl08|dressed_sharp|-0.7707|0.324|0.676|0.0|"RT @dressed_sharp: There s nothing patriotic about accepting a fraudulent election, real Americans will go to court if #trump loses because"
DadandBuried|dadandburied|-0.5719|0.171|0.829|0.0|"""What Trump is really doing is legitimizing hate for a large segment of the population that has a lot of it.""https://t.co/yfQwbMxHXg"
zanesholtz|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
sw7617|Henryyearwood1|-0.6124|0.25|0.75|0.0|RT @Henryyearwood1: @Serenity_Seas @FedUp137 @JackPosobiec of course the hacks will no worries West Florida will vote Trump
nickiloc|GaryLineker|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
nickiloc|twitter|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
Txndras_|SheHatesJacoby|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
Txndras_|twitter|0.0|0.0|1.0|0.0|RT @SheHatesJacoby: President Obama still roasting Trump.. 4th Quarter Obama been shooting 100%  https://t.co/xGBnJVL5Lu
wbcurley|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
wbcurley|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
justquincy_|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
justquincy_|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
tamaraleighllc|DonaldJTrumpJr|0.4753|0.0|0.866|0.134|RT @DonaldJTrumpJr: FOX NEWS EXIT POLL: 87% of voters believe my father is the true change candidate. #MAGA GO VOTE! #TRUMP
Brianna13Ortiz|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
rosado_jm|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
lesliegtz_|fuckowiak|0.3182|0.0|0.85|0.15|"RT @fuckowiak: please remember to vote, unless you're voting for trump then stay home"
kmsangelica|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
kmsangelica|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Barnett_59|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
ViciousVeeeeeee|flawedfacade|0.0|0.0|1.0|0.0|RT @flawedfacade: Y'all talmbout a Trump presidency turning the clock back 500 years when in reality it'll turn the clock back less than 50
Cuffs_No_Hoes|TheHomieLos|0.0|0.0|1.0|0.0|"RT @TheHomieLos: ""Vote for Hillary to keep Trump out of office""...I get it. But I need way more than that homie."
ReconmomC|RapinBill|0.8349|0.0|0.745|0.255|"RT @RapinBill: Numbers were looking good, now they are looking Great for Trump! Keep it up! Get Everybody you can To Vote for Trump! #Elect"
209twitch|MaxMeleganich|-0.1531|0.348|0.652|0.0|@MaxMeleganich @inshaIlah awkward https://t.co/4vRGCllGBU
209twitch|nytimes|-0.1531|0.348|0.652|0.0|@MaxMeleganich @inshaIlah awkward https://t.co/4vRGCllGBU
BrandonMPuleo|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
BrandonMPuleo|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
drginareghetti|fanofcars|-0.3432|0.124|0.876|0.0|RT @fanofcars: #Trump#FBIDirector #CNN#voterfraud Who takes this seriously? How are these corrected b4 Nov 8th? Who is responsible?W
LULUBELLE1000|FaithRubPol|0.6705|0.0|0.814|0.186|"RT @FaithRubPol: It is impossible for Trump to #maga because he will give up our values. As Lincoln said, ""let us have faith that RIGHT mak"
melsmonts|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
developertest09|twitter|0.0|0.0|1.0|0.0|Ouch for Hillary. Even if Indies only break for Trump +5% it would be OUCH. https://t.co/RqBOillxUd
AndrewsCosta4|IBTimes|-0.4939|0.225|0.775|0.0|RT @IBTimes: Mosques across the country are fearful heading into #ElectionNight https://t.co/5YcGl0CFPS
AndrewsCosta4|ibtimes|-0.4939|0.225|0.775|0.0|RT @IBTimes: Mosques across the country are fearful heading into #ElectionNight https://t.co/5YcGl0CFPS
phoebe__warren|KayBurley|0.0|0.0|1.0|0.0|RT @KayBurley: BREAK: George W Bush and wife Laura say they didn't vote for Trump #Election2016
guwop_07|Iplayforthefun|0.3818|0.0|0.88|0.12|RT @Iplayforthefun: I just thought about Donald trump becoming president and I calmed myself down by remembering j. Cole when double platin
_adornk|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_adornk|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
danialx|Sporf|-0.3182|0.173|0.827|0.0|RT @Sporf: BREAKING: Stone Cold interrupts the Donald Trump rally.  #ElectionDay( @thrillis4)https://t.co/zJZAmoHlNY
danialx|twitter|-0.3182|0.173|0.827|0.0|RT @Sporf: BREAKING: Stone Cold interrupts the Donald Trump rally.  #ElectionDay( @thrillis4)https://t.co/zJZAmoHlNY
worldnews_net|abcnews|0.0|0.0|1.0|0.0|How Donald Trump Is Spending Election Night https://t.co/zmNZ6HvF1w #abcnews #abc #news
DavidMk11|Fatality_89|0.0|0.0|1.0|0.0|RT @Fatality_89: Trump Cake https://t.co/UIIioGmnXr
DavidMk11|twitter|0.0|0.0|1.0|0.0|RT @Fatality_89: Trump Cake https://t.co/UIIioGmnXr
lgbtqtyIer|ridevocals|-0.4588|0.146|0.778|0.075|"RT @ridevocals: WHY ARE PEOPLE VOTING TRUMP BECAUSE ""HILLARY IS A CRIMINAL"" WHEN THE FBI ALREADY CLEARED HER AND TRUMP IS GOING TO COURT FO"
sms442|DanScavino|0.0|0.0|1.0|0.0|RT @DanScavino: Trump Campaign Headquarters-'TOP CANDIDATE QUALITY: CAN BRING CHANGE:TRUMP: 82%CLINTON: 13%#iVoted #ElectionNight #MAGA
buckeyery|TattooedNnerdy|0.0|0.0|1.0|0.0|RT @TattooedNnerdy: #voted @TYTNetwork @HillaryClinton @realDonaldTrump #ElectionNight Hillary+Trump=  https://t.co/1BwijJ7flw
buckeyery|twitter|0.0|0.0|1.0|0.0|RT @TattooedNnerdy: #voted @TYTNetwork @HillaryClinton @realDonaldTrump #ElectionNight Hillary+Trump=  https://t.co/1BwijJ7flw
TYMZUS666|KayzoMusic|0.4215|0.0|0.714|0.286|RT @KayzoMusic: Do u think Donald trump likes riddim
king23tahj|kilhoes|0.6597|0.0|0.649|0.351|"RT @kilhoes: ""Do you think Trump has a chance of winning""  #ElectionNight https://t.co/bV9oRNHTVR"
king23tahj|vine|0.6597|0.0|0.649|0.351|"RT @kilhoes: ""Do you think Trump has a chance of winning""  #ElectionNight https://t.co/bV9oRNHTVR"
ymirius|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
ymirius|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
GuruVShetty|madhukishore|0.3612|0.0|0.848|0.152|RT @madhukishore: Like for Hillary or Retweet for Trump #ElectionDay #ElectionNight #ElectionFinalThoughts #USElection2016 #USADecides #Vot
drewjacorey_|Iam_Kinnaird|0.3818|0.122|0.667|0.211|RT @Iam_Kinnaird: It was a no brainer that Trump was gonna win Indiana and Kentucky..
AmyJoyHagen|blahblah8976|0.0|0.0|1.0|0.0|@blahblah8976 @MotherJones oh I did vote!!! For trump! #trumptrain #womenfortrump #michiganfortrump
Rayneeebow|gvbigz|-0.5795|0.178|0.822|0.0|"RT @gvbigz: no, we rly can't be friends if u cast your vote for Trump not understanding the implications exceed that of simply holding ""dif"
IlinaMilada|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
IlinaMilada|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ZhukovElmar|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ZhukovElmar|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
GOPbattle2016|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
SlaaayTf|_AsToldByShayy_|0.7488|0.101|0.629|0.27|RT @_AsToldByShayy_: If Donald trump wins !!! Let's all not go to work tomorrow and scare the shit out of the government  #Retweet
mikemyres12|AlGaldi|0.0|0.0|1.0|0.0|"RT @AlGaldi: #PresidentialElection sports comps.  I have #Trump as Steinbrenner, #Hillary as #ARod &amp; the race as a whole as the #MalaceAtTh"
alicezinawhitt|TheHazelHayes|0.0|0.0|1.0|0.0|"RT @TheHazelHayes: #Trump is a big, fat, orange, Putin-loving, gay-bashing, hate-mongering, wall-building, gun-toting, wig-wearing, pussy-g"
JosieNano|twitter|0.0|0.0|1.0|0.0|Call trump hotline and report them !!!!!! https://t.co/0OFTJYAuNJ
patriot1cavalry|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
patriot1cavalry|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
alabaluu|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
alabaluu|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
Satch7Eddie|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
Ellojoe|chrislhayes|0.0|0.0|1.0|0.0|"RT @chrislhayes: After waiting until almost *literally* the last moment, Toomey votes and says he voted for Trump."
gaidargorbuno10|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
gaidargorbuno10|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
worldnews_net|latimes|0.0|0.0|1.0|0.0|Former President George W. Bush didn't vote for Donald Trump https://t.co/1CVbfh9MRJ #LosAngelesTimes #latimes #news
VJ_Ostrowski|twitter|-0.3621|0.174|0.711|0.115|"Trump: ""this was very VERY unfair to me. Many of my supporters are gamer weaboos. They stayed home now."" https://t.co/7u7PvI1xWW"
LuckymeEva|h1llary4prez|0.4019|0.0|0.876|0.124|RT @h1llary4prez: #ImWithHer because she can work with both parties. Trump has proven he can work with neither. #Election2016 #ElectionDay
irishsox3|scottzolak|0.0|0.0|1.0|0.0|@scottzolak @Dan_Shaughnessy @BostonGlobe shut up shank. Go Trump!
WhosGoneGalt|GiveMeLibertyUS|0.4939|0.0|0.878|0.122|"RT @GiveMeLibertyUS: Come on late voters in FL, PA, Ohio, etc.  Get out and vote 4 Trump - let's seal the Deal.  Let's save America - Make"
miraculashton|HillaryClinton|-0.743|0.249|0.751|0.0|"RT @HillaryClinton: ""If you believe that racism and sexism and bigotry have no place in our country...you need to vote."" https://t.co/nIOvu"
miraculashton|t|-0.743|0.249|0.751|0.0|"RT @HillaryClinton: ""If you believe that racism and sexism and bigotry have no place in our country...you need to vote."" https://t.co/nIOvu"
amandahoopes|CNN|0.0|0.0|1.0|0.0|"RT @CNN: Trump: We're going to build a wall. Who's paying for it?Crowd: ""Mexico""Trump: ""100 percent"" https://t.co/HEdS8bVcgo"
amandahoopes|twitter|0.0|0.0|1.0|0.0|"RT @CNN: Trump: We're going to build a wall. Who's paying for it?Crowd: ""Mexico""Trump: ""100 percent"" https://t.co/HEdS8bVcgo"
Trumppatriot2|KellePsychic|0.8176|0.0|0.653|0.347|RT @KellePsychic: Trump voters and nation lots of positive energy around him have faith our prayers have manifested.#TrumpPence16 @DonaldTr
taliadelrey|THOTJAI|0.5719|0.0|0.821|0.179|RT @THOTJAI: if donald trump wins the election I will paypal 100 dollars to everyone that retweets this #ElectionDay
ALESSSANDROPERU|DanScavino|0.5473|0.0|0.757|0.243|@DanScavino @TeamTrump @mike_pence @Trump @atvmasnoticias @RPPNoticias @cala  ***CONGRATULATIONS***NEW PRESIDENT UNITED STATES ***TRUMP***
patriciamcivor1|rooshv|0.4215|0.0|0.833|0.167|"RT @rooshv: My mother, sister, father, and brother all voted for Trump. Bless them. https://t.co/ivfqIuAKbD"
patriciamcivor1|twitter|0.4215|0.0|0.833|0.167|"RT @rooshv: My mother, sister, father, and brother all voted for Trump. Bless them. https://t.co/ivfqIuAKbD"
Patmijares_|salazaroreste61|0.2516|0.076|0.807|0.117|"RT @salazaroreste61: All my co-workers are Trump supporters, needless to say it's very awkward being the only Hispanic (Mexican to be speci"
KimberMolyneux|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
KimberMolyneux|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
holcomb_todd|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you voted for TRUMP! #ElectionDay #Vote #Vote2016
MpressT|jorgeramosnews|-0.4215|0.149|0.851|0.0|RT @jorgeramosnews: Univision's Jorge Ramos says Trump's snub of Latino media will cost him https://t.co/bZOuqjoLKE via @CNNMoney
MpressT|money|-0.4215|0.149|0.851|0.0|RT @jorgeramosnews: Univision's Jorge Ramos says Trump's snub of Latino media will cost him https://t.co/bZOuqjoLKE via @CNNMoney
stevenj60329854|QualityStrange|-0.6369|0.245|0.755|0.0|RT @QualityStrange: @rj47972891 This is a fake poll making the rounds to get Trump voters to stay home. Disregard
Mahoney2John|vivelafra|0.0|0.0|1.0|0.0|@vivelafra trump trump president
davidpwil|MissLizzyNJ|0.0|0.0|1.0|0.0|"RT @MissLizzyNJ: Remember, Hillary will take an early lead in exit polls which will change drastically, once Trump voters get out of work."
KramerFry|Swordsmanx10|0.5719|0.0|0.812|0.188|"RT @Swordsmanx10: WIKILEAKS 1-35 BREAKING NEWS: Donald Trump Wins Florida, OH, NC Despite ... https://t.co/s8Kw4VjCVX via @YouTube"
KramerFry|youtube|0.5719|0.0|0.812|0.188|"RT @Swordsmanx10: WIKILEAKS 1-35 BREAKING NEWS: Donald Trump Wins Florida, OH, NC Despite ... https://t.co/s8Kw4VjCVX via @YouTube"
gnarruto|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Dj2Brazy|dvpecain|0.3094|0.086|0.774|0.14|"RT @dvpecain: 2016- Trump won't win2017- President Trump can't do that , can he?2018- say u watching the hunger games tonight? I hope m"
thewickedlilith|CurveMe|0.6633|0.0|0.772|0.228|RT @CurveMe: IF TRUMP WINS THE ELECTION   IM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICAGOODMORNINGSAN DIEGO
GoykhmanAlla|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: Trump now leading IN by 45 points.  RCP has him by 10.  Something is happening.
RebeccaGrant77|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
RebeccaGrant77|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
jujuuballs|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
jujuuballs|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
JustAcceptFate|NBCNewYork|0.0|0.0|1.0|0.0|@NBCNewYork D Trump shall conquer clinton
Gfabgab|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Gfabgab|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
svogel2|RichardGrenell|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
svogel2|twitter|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
geraldin_oe|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
DemiIsAll|ddlsbodysay|0.4995|0.0|0.773|0.227|RT @ddlsbodysay: RT for Demi Lovato LIKE for Donald Trump #ElectionDay https://t.co/0olnXz8Dcg
DemiIsAll|twitter|0.4995|0.0|0.773|0.227|RT @ddlsbodysay: RT for Demi Lovato LIKE for Donald Trump #ElectionDay https://t.co/0olnXz8Dcg
thelilkait|frandmnd|0.7003|0.0|0.547|0.453|RT @frandmnd: Good morning to everyone except trump supporters
willluv1Dalways|twitter|0.6996|0.186|0.319|0.494|Pretty much! I hope the racists Trump supporters don't win:) https://t.co/AT414dUNIW
ncisissick|270towin|0.0|0.0|1.0|0.0|"This is what I think will happen tonight. However, Trump could flip a few other blue states, such as; Nevada,... https://t.co/fCXXUjbQYU"
TrumpAmerica17|michaeljohns|0.0|0.0|1.0|0.0|"RT @michaeljohns: #Florida: If you are in line by 7pm ET tonight, you can still vote. 20 minutes:#TeaParty #Trump2016 #TrumpTrain #Trum"
Smokey91199|szeachmoment|0.0772|0.0|0.885|0.115|RT @szeachmoment: @theglobaluniter @DonaldJTrumpJr panhandle dweller here. Everyone I know voted Trump.
MadameRamotswe|karlazabs|-0.5106|0.171|0.829|0.0|Meet The Abused Workers Who Sewed Donald Trump Clothing For A Few Dollars A Day https://t.co/jJ28Li8JrJ via @karlazabs @buzzfeednews
MadameRamotswe|buzzfeed|-0.5106|0.171|0.829|0.0|Meet The Abused Workers Who Sewed Donald Trump Clothing For A Few Dollars A Day https://t.co/jJ28Li8JrJ via @karlazabs @buzzfeednews
janakatharine8|twitter|0.6249|0.0|0.806|0.194|Make America Great Again hats bookend the stage inside the Hilton ballroom for Donald Trump's #ElectionNight event https://t.co/eKSizUA3og
MrsLeeJooheon|trblheaux|0.5719|0.0|0.778|0.222|RT @trblheaux: We need to plan a twitter meetup at the plantation when Trump wins
TrippyyTayy|FunniestVines|0.6408|0.0|0.68|0.32|RT @FunniestVines: This guy electrified his Trump sign LMFAO  https://t.co/uXwAXer6PC
TrippyyTayy|twitter|0.6408|0.0|0.68|0.32|RT @FunniestVines: This guy electrified his Trump sign LMFAO  https://t.co/uXwAXer6PC
doparrish51|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
doparrish51|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
J0HN_chambers|lmNotWhite|0.5106|0.093|0.662|0.245|RT @lmNotWhite: If Trump wins I'll pay everyone $5 who RTs this.
yarike|vandives|0.4753|0.0|0.853|0.147|"RT @vandives: I just voted for our next president, Donald J. Trump  a true American patriot &amp; the ultimate MADMAN!#MAGA3X #MAGASELFIE "
itmealexx|DonaldJTrumpJr|0.5696|0.0|0.872|0.128|"RT @DonaldJTrumpJr: If you have friends in MI, OH, FL, PA -- CALL THEM and tell them to VOTE TRUMP! You can make a difference! #MAGA #Tru"
eightzenuff|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
s0phicee|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
s0phicee|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
asperry3|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
helenecdexter|GaryLineker|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
helenecdexter|twitter|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
jaira13s|FranchiseRocks|-0.9195|0.547|0.453|0.0|RT @FranchiseRocks: Damn bro. Hillary and Trump are the fucking devil. We're fucked.
_Smeg|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
_Smeg|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
RealVinnieJames|Ekatherene|0.34|0.0|0.769|0.231|@Ekatherene @Always_Trump Games people play. Deleting it now. -VJ
MuttonMusic|Cain_Unable|0.0|0.0|1.0|0.0|"RT @Cain_Unable: I just tried to Vote Trump &amp; the staff wouldn't let me just because I'm ""in Kent"" &amp; ""this is a Tesco self service checkout"
DADIG123|markcritch|0.0|0.0|1.0|0.0|RT @markcritch: I assume this was because #Trump had never voted before and didn't know how #ElectionDay https://t.co/wdzWvjKGLH
DADIG123|twitter|0.0|0.0|1.0|0.0|RT @markcritch: I assume this was because #Trump had never voted before and didn't know how #ElectionDay https://t.co/wdzWvjKGLH
mamasaurusof2|thehill|0.4019|0.0|0.863|0.137|RT @thehill: Twitter users speculate: Is Cindy McCain's white pant suit a show of support for Clinton? https://t.co/ALR17pjOX1 https://t.co
mamasaurusof2|thehill|0.4019|0.0|0.863|0.137|RT @thehill: Twitter users speculate: Is Cindy McCain's white pant suit a show of support for Clinton? https://t.co/ALR17pjOX1 https://t.co
0321jail|MightyBusterBro|0.0|0.0|1.0|0.0|RT @MightyBusterBro: .A MUST SEE VIDEOINSPIRATIONAL MOMENTFINAL TRUMP RALLY@realDonaldTrump#VOTE  #ElectionDay #MyVote2016 #MAGA htt
gehenna1888|ananavarro|-0.2732|0.087|0.913|0.0|"RT @ananavarro: Hey Nevadans, u know why Trump is suing? To keep Hispanics from polls b/c he knows we're voting against him. Redouble your"
xjenncarv|_carolineotoole|0.6597|0.0|0.787|0.213|"RT @_carolineotoole: If you vote Trump tomorrow, make sure explain to your gay, trans, female, black, Latina/o, and Muslim friends why they"
9ERSorBUST|YouTube|0.0|0.0|1.0|0.0|"Scientific Poll Shows Trump With ""Yuge"" Lead in Swing States https://t.co/WmQIJ3Ex0H via @YouTube"
9ERSorBUST|linkis|0.0|0.0|1.0|0.0|"Scientific Poll Shows Trump With ""Yuge"" Lead in Swing States https://t.co/WmQIJ3Ex0H via @YouTube"
6nsinvt|chicoscperez|-0.4019|0.144|0.856|0.0|"RT @chicoscperez: Donald Trump Has a Millennial Problem, and It Could Reshape American Politics via @thenation https://t.co/B12LXlu0Xf #TNT"
6nsinvt|linkis|-0.4019|0.144|0.856|0.0|"RT @chicoscperez: Donald Trump Has a Millennial Problem, and It Could Reshape American Politics via @thenation https://t.co/B12LXlu0Xf #TNT"
izzyfizzy1123|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
izzyfizzy1123|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
BIGMONEYMETTA|BuzzFeedNews|0.5859|0.0|0.853|0.147|RT @BuzzFeedNews: Here we go: Kentucky is one of the first polls to close and BuzzFeed News expects Donald Trump to win  https://t.co/OMYv
BIGMONEYMETTA|t|0.5859|0.0|0.853|0.147|RT @BuzzFeedNews: Here we go: Kentucky is one of the first polls to close and BuzzFeed News expects Donald Trump to win  https://t.co/OMYv
Kare_FreeTrudy|9EtherKing|-0.6359|0.224|0.776|0.0|@9EtherKing by the looks of it Trump leading so wrong question . Question is wah time the boat leave to Africa ?
GreggBeratan|UniteWomenWV|-0.1982|0.161|0.646|0.193|RT @UniteWomenWV: Please share this article on why @realDonaldTrump is so dangerous for people w/ disabilities! #CripTheVote @bustle https:
CamillaSposito|DrPresidentPat|-0.8208|0.274|0.726|0.0|RT @DrPresidentPat: DONALD TRUMP'S SON MAY HAVE JUST DISQUALIFIED HIS VOTE FOR HIS OWN FATHER I CANNOT BREATHE IMAGINE BEING THIS DUMB http
HotdesertAz65|Judgenap|-0.3544|0.125|0.794|0.08|@Judgenap VOTE TRUMP AND A NEW GOVT THAT WILL DO THE RIGHT THING AND NOT ALLOW ANYONE TO LIVE ABOVE THE LAW !!! NO ONE IS ABOVE THE LAW !
JohnburW|youtube|0.5754|0.0|0.682|0.318|BLACKS AND LATINOS STARTING TO SUPPORT DONALD TRUMP! https://t.co/ihiwTW1fh5
josephiykech|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
ahbying|politico|-0.0191|0.107|0.893|0.0|Tom Brady's wife says the QB isn't backing Trump https://t.co/ensM9rAJk0
Mitchllryancain|Atom_Murray|0.2263|0.0|0.863|0.137|RT @Atom_Murray: Okay. Now I'm done with the Trump Cake tweets. #ElectionNight https://t.co/4jtsTFA9PR
Mitchllryancain|twitter|0.2263|0.0|0.863|0.137|RT @Atom_Murray: Okay. Now I'm done with the Trump Cake tweets. #ElectionNight https://t.co/4jtsTFA9PR
PhatLikeBuddha|twitter|-0.3818|0.191|0.809|0.0|This the final boss fight for anyone tryna vote against Trump https://t.co/7C4kB9Ii44
MattPosorske|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
Sauje|damaninthearena|0.0|0.0|1.0|0.0|RT @damaninthearena: @Vendetta92429 @antimarxis_ this map is BS!! I'm in southern Cali and in a line of 50+ people; Black White Hispanic As
fangpusskins|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
fangpusskins|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
nrsMichigan|RichardGrenell|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
nrsMichigan|twitter|0.7425|0.089|0.567|0.344|RT @RichardGrenell: Completely true. The LGBT community is supporting Trump like no other GOP presidential candidate before. https://t.co/M
smaragdkolesni2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
smaragdkolesni2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
Wordsmiter|Miami4Trump|0.7003|0.0|0.766|0.234|RT @Miami4Trump: Trump Cares About Inner Cities And Improving Education. He's discussed This For Over 30 YEARS #VoteTrump He Will #MAGA#El
LeeLee_Ri|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
LeeLee_Ri|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
PatriciaArnona|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you voted for TRUMP! #ElectionDay #Vote #Vote2016
3rdwheelawkward|RealTimers|0.1027|0.082|0.82|0.098|"RT @RealTimers: ""Anybody sitting on the sidelines right now or deciding to engage in a protest vote that's a vote for Trump.""  @POTUS #U"
ShelleyOberg|EricTrump|0.0|0.0|1.0|0.0|@EricTrump @realDonaldTrump go trump #draintheswamp
davidappell|kurteichenwald|0.0516|0.093|0.806|0.101|"RT @kurteichenwald: Ive been asked several times what happens if Trump loses &amp; won't concede. The answer is: Nothing. It's a courtesy, not"
heatherxstarrr|polaroidbones|-0.607|0.184|0.816|0.0|RT @polaroidbones: DONT SPLIT THE DEMOCRATIC VOTE TOMORROW CAUSE YOU DONT WANNA BE STUCK HILLARY OR TRUMP! ITS ONLY GONNA LEAVE US WITH TRU
abern918|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
Leeceea1|Trump2016News|0.0|0.0|1.0|0.0|"RT @Trump2016News: Republicans: I know you're all busy WORKING, but don't put off voting at 5PM! Trump never gave up on you; don't give up"
conciousIy|troyesivan|-0.3182|0.133|0.867|0.0|RT @troyesivan: i dont mean to be a tease but....like...imagine not having to hear about donald trump anymore 
Horsies_MUT|Dona1dTrumpMUT|-0.3182|0.187|0.813|0.0|@Dona1dTrumpMUT so do you stay with the same @ if Trump loses?
moneeyy___|StahrMilan|-0.658|0.16|0.84|0.0|RT @StahrMilan: And to see people still down talking Hillary! Shut up bitch! When Bernie was running YALL ain't vote now it's Hillary and t
TheSteeldawn|Khaixur|-0.743|0.259|0.741|0.0|"@Khaixur If it's proven that clinton rigged states with voter fraud and election rigs, then trump ends up being right."
DrMorien1|mitchellvii|0.5719|0.0|0.85|0.15|"RT @mitchellvii: Romney won Brevard County by 36,000 votes in 2012.  I calculate Trump leads it by 52,000 votes.  +16,000 votes for Trump o"
hector_bolt|mrmichaelpersad|-0.7233|0.252|0.652|0.096|"RT @mrmichaelpersad: [obama running]""WHAT RELIGION IS HE?? WHERE WAS HE BORN!?! HES A TERRORIST"" [trump running]""dont act like you ne"
AMLx3|simplysydd|-0.8768|0.339|0.587|0.073|RT @simplysydd: I dead ass I know ppl that voted for Donald trump. Like ppl I was close to. Ppl really are closeted racists and you don't e
SaBrown93|MicaBurton|0.4019|0.218|0.489|0.293|@MicaBurton i hope for your countries sake Hillary wins. no country should be burdened with Trump
taehyungstounge|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
LGarchomp|RobZyo|0.372|0.075|0.791|0.134|RT @RobZyo: 2016: Trump won't win2017: President Trump can't do that can he?!2018: So you watching the Hunger Games tonight? I hope my di
lyn_gb|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
lyn_gb|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
ConservativLuke|Guy75356686|-0.5423|0.241|0.759|0.0|RT @Guy75356686: @mflynnJR @mitchellvii we are voting our ass off for Trump
pteacherinme|seethew0rld|0.0|0.0|1.0|0.0|RT @seethew0rld: #FL #PCB Panhandle GET OUT THE VOTE #Trump https://t.co/VygXKMIuSC
pteacherinme|twitter|0.0|0.0|1.0|0.0|RT @seethew0rld: #FL #PCB Panhandle GET OUT THE VOTE #Trump https://t.co/VygXKMIuSC
stevengale57|pudcast245|0.7003|0.0|0.756|0.244|RT @pudcast245: I give it about 4-5 hrs before the #deplorable #Trump supporters with #Pepe profiles start disappearing from Twitter. Good
skywolfangel|DilaChuu|0.3612|0.0|0.706|0.294|RT @DilaChuu: Not to say I like trump
lavrentevaminn2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
lavrentevaminn2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
memeswearmatty|letters2donald|0.3612|0.0|0.865|0.135|"RT @letters2donald: Children's letters to Donald Trump:  Does Melania like you cause shes a lier too?April H., age 8"
blancaportill21|soul4ever|-0.3818|0.167|0.833|0.0|"RT @soul4ever: Trump is rude and unsophisticated, he disrespects anyone but himself. I can't believe how many people vote for him.#Election"
JR777771|kindcutesteve|-0.4404|0.153|0.847|0.0|RT @kindcutesteve: Latino Voter Wall Will Block Trumps Path to White House (thank you Latino's)#p2 #TNTweeters #USLatinohttps://t.co/q2P
JoshuaMLopez_|twitter|0.5994|0.138|0.545|0.316|"Suuuuure, buddy. Everything's a fraud with you people. Grow up and accept that Donald Trump has a pretty good chanc https://t.co/OPi8GiUrEO"
hyejenog|aeriaIview|0.3612|0.0|0.872|0.128|@aeriaIview theres a guy named Bolsonaro he's like trump but.. worse(?) and he's thinking about becoming a president in 2018
JoLoDiBenedetto|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
reisegrrl1|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
Nhevi_XO|theyearofelan|-0.6566|0.196|0.804|0.0|RT @theyearofelan: Wouldn't it be amazing if Trump lost New York by one vote because his son illegally took a photo of his completed ballot
donah1121|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: VOTER FRAUDVotes flipped from Trump to Clinton in Pennsylvania.#ElectionDay #Voted #Vote2016 https://t.co/EKy4TqxTiX
donah1121|twitter|0.0|0.0|1.0|0.0|RT @America_1st_: VOTER FRAUDVotes flipped from Trump to Clinton in Pennsylvania.#ElectionDay #Voted #Vote2016 https://t.co/EKy4TqxTiX
carolineeileen_|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
carolineeileen_|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
UrbanismAvenger|ajplus|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
UrbanismAvenger|twitter|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
jurrjurrtbull|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
carbidethung|mitchellvii|0.7998|0.0|0.736|0.264|RT @mitchellvii: The last RCP Poll had Trump winning KY by 17.  He is currently winning by 52 points.Monster vote?  Dem crossovers?
williamcreedcox|vitweet|0.0|0.0|1.0|0.0|MN Voters We Need Your VotesPlease don't do anything after work except VOTE TRUMP! Get to your  #DrainTheSwamp https://t.co/aHVAa5Dccp
CHRISTINA2A12|mrbeercrusher|0.0|0.0|1.0|0.0|RT @mrbeercrusher: Expect a Trump victory in North Carolina announced around eight o'clock eastern time. Trump up 3.7% in the average of ex
MrEdTrain|surfermom77|0.0|0.0|1.0|0.0|"RT @surfermom77: Twitter &amp; FB R begin inundated wt reports of Elec.fraud, voting irregularities &amp; discrimination against Trump Votershttps"
USA_with_Trump|NAAlmodovar|0.0|0.0|1.0|0.0|RT @NAAlmodovar: All I hear is how crooked H is as I wait on line in small town Idaho. Line is over 60 minutes long.
BrandConverts|costareports|0.0|0.0|1.0|0.0|"RT @costareports: On the phone w/ Giuliani. He just left Trump's apt. Said Trump is ""watching everything even tho I'm telling him not to."""
SWFCStefan|GaryLineker|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
SWFCStefan|twitter|0.6808|0.0|0.741|0.259|RT @GaryLineker: I must say your ability to continually tweet from deep inside Trump's bowels is rather impressive. https://t.co/eBgeY3Nell
IRepBlakkk|TheOiz|0.7964|0.0|0.712|0.288|"RT @TheOiz: In the event Donald Trump wins, I'm just hoping people of color can get a day off of work/school/everything for emotional distr"
Mr3lsewhere|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
Mr3lsewhere|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
tony_ganzer|NickCastele|0.0|0.0|1.0|0.0|RT @NickCastele: Director of @cuyahogaboe says rumored self-appointed Trump election observers didn't show up at polling places here.
HiKambrya|Deadspin|0.0|0.0|1.0|0.0|RT @Deadspin: The Trump campaign wants to make names of Nevada poll workers public. Judge's response: https://t.co/tes99IMbbH
HiKambrya|twitter|0.0|0.0|1.0|0.0|RT @Deadspin: The Trump campaign wants to make names of Nevada poll workers public. Judge's response: https://t.co/tes99IMbbH
MADE__USA|09BRAININJURY|0.6523|0.0|0.75|0.25|RT @09BRAININJURY: @deplorablelori MY WIFE AND I VOTED FOR MY HERO AND IDOL MR.TRUMP TONIGHT
Tyreke_p|NathanZed|0.5719|0.0|0.866|0.134|RT @NathanZed: if trump wins im moving to my grandmas house. she still live in america this don't got anything to do with politics I just m
halebopp_79|tinnnies|0.3182|0.09|0.748|0.162|RT @tinnnies: I'm scared to wake up tomorrow and see that trump has won it will be the same heart breaking feeling as waking up to brexit
lilrascal01|iResistAll|0.6249|0.0|0.779|0.221|"RT @iResistAll: BREAKING: Durham County, NC to extend voting in Democrat areas because Trump is winning the state. #electionday #ElectionN"
nickstuart118|64_bit_hero|0.0|0.0|1.0|0.0|RT @64_bit_hero: Donald Trump sticks PS1 memory cards up his arse
goldnbeak|jaketapper|0.3566|0.0|0.894|0.106|"RT @jaketapper: But then Trump couldn't run, since his mom and paternal grandparents weren't born in the US. So, um, yeah. https://t.co/7Ux"
goldnbeak|t|0.3566|0.0|0.894|0.106|"RT @jaketapper: But then Trump couldn't run, since his mom and paternal grandparents weren't born in the US. So, um, yeah. https://t.co/7Ux"
BlastingNews|us|0.0|0.0|1.0|0.0|#election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR https://t.co/AfJAdNdbSU
ssammysuave|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
Avocadohomo|lntroset|0.8969|0.0|0.67|0.33|RT @lntroset: Today is Election Day so I thought I would share the loving someone lyrics with you guys bc this world needs more love and le
allison_fether|chelseahandler|0.3612|0.0|0.906|0.094|"RT @chelseahandler: Stevie Wonder said that voting for Trump is like asking me to drive."" Id rather have Stevie as my Uber driver than Tr"
feeIthebreeze|twitter|0.6239|0.0|0.631|0.369|"""And the winner is Donald Trump!"" #ElectionNight https://t.co/7lxTTjXGYu"
jakeroberts2015|YahooNews|-0.8689|0.353|0.647|0.0|RT @YahooNews: WATCH LIVE: GOP pollster @FrankLuntz says Its a vote between a liar and a lunatic &amp; people will choose the liar https://t
jakeroberts2015||-0.8689|0.353|0.647|0.0|RT @YahooNews: WATCH LIVE: GOP pollster @FrankLuntz says Its a vote between a liar and a lunatic &amp; people will choose the liar https://t
bmelton00|UntamedJeaux|-0.25|0.104|0.833|0.063|RT @UntamedJeaux: Illegals complain about trump wanting to deport them.. Go through the legal process to become a fucking citizen of the U.
AaronSims31|March_for_Trump|-0.5766|0.186|0.74|0.074|RT @March_for_Trump: An urgent message on #Voterfraud coming from @cubans4trump. REPORT VOTER FRAUD: 855 976 1200 (Trump Lawyer Team).; #El
GaryAddington|_Makada_|-0.2714|0.185|0.694|0.121|RT @_Makada_: REPORT: Man Attacks Female Trump Supporter at Florida Polling Station! #ElectionDay https://t.co/Zw4MbGuxvP
GaryAddington|thegatewaypundit|-0.2714|0.185|0.694|0.121|RT @_Makada_: REPORT: Man Attacks Female Trump Supporter at Florida Polling Station! #ElectionDay https://t.co/Zw4MbGuxvP
JimenezValejm27|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
JimenezValejm27|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
perrya11|DonaldJTrumpJr|0.7906|0.0|0.75|0.25|RT @DonaldJTrumpJr: FINAL PUSH!Lets RT THIS TO A TRUMP VICTORY!RT if you want to see TRUMP WIN TONIGHT! #MAGA Not too late to vote! G
Chitown1216|MattGertz|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
Chitown1216|twitter|-0.7269|0.337|0.663|0.0|RT @MattGertz: CNN's Jake Tapper: Trump is lying about nationwide voting machine problems. https://t.co/HfPt0wHxmp
shayne571|twitter|-0.4019|0.172|0.828|0.0|Main problem with Republicans. Still think Clinton was beatable by someone Trump beat. https://t.co/vrbxb1xRqf
Javi_GV_ATM|mrbeercrusher|-0.7672|0.259|0.741|0.0|RT @mrbeercrusher: #ElectionDay SHOCK Exit Polls have Clinton campaign in panic mode:Trump up 3.4% in PATrump up 2.1% in MichTrump up 3
kimlitwicki|TeamTrump|0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
kimlitwicki||0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
princejaygt|UglyGod|-0.5106|0.121|0.879|0.0|RT @UglyGod: It means yall shoulda fuckin listened &amp; kept Bernie Sanders as an option cause now we all look dumb af choosing between Hillar
therightworks|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
therightworks|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
asiyakondratev2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
asiyakondratev2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
cliffordtopham|WDFx2EU8|0.0|0.0|1.0|0.0|RT @WDFx2EU8: BREAKING: TRUMP is getting 27% of latino vote based on early exit vote. Overperforming projections https://t.co/PJvl40rsFM
cliffordtopham|twitter|0.0|0.0|1.0|0.0|RT @WDFx2EU8: BREAKING: TRUMP is getting 27% of latino vote based on early exit vote. Overperforming projections https://t.co/PJvl40rsFM
UKolizer|uk|0.0|0.0|1.0|0.0|George Bush did not vote for Donald Trump https://t.co/JuQRXrEK3C https://t.co/DP0Nq8oIQf
constantino_sam|pinterest|-0.8208|0.457|0.543|0.0|TRUMP THAT BITCH - ANTI HILLARY PRO TRUMP POLITICAL BUMPER STICKER https://t.co/hlE23UztMY
Nina_mk_|AmandaMiIIs|-0.4404|0.266|0.734|0.0|RT @AmandaMiIIs: If you're voting for trump block me
Savannah_JeaD|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
Savannah_JeaD|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
britneygarcia_|ari_brendan|0.4939|0.072|0.72|0.208|RT @ari_brendan: @HuskJonathan alright Jonny seriously enough with the ignorance.Lets just hope America is still up and running if inhumane
dronerecovery|neko_designer|0.3182|0.0|0.839|0.161|"@neko_designer @ShimermanArmin ""please see the treatment of trump"" Appeal to hypocrisy, second count."
tifmcclure|mitchellvii|0.7998|0.0|0.736|0.264|RT @mitchellvii: The last RCP Poll had Trump winning KY by 17.  He is currently winning by 52 points.Monster vote?  Dem crossovers?
Piercepierce87|BetteMidler|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
Piercepierce87|twitter|-0.5852|0.256|0.744|0.0|RT @BetteMidler: I guess the Trump men don't really trust their wives!!! https://t.co/E2Vyz2V0fp
_PurpleUnicorns|l4444k|0.0|0.0|1.0|0.0|RT @l4444k: Snoop Dogg @ Donald Trump Roast https://t.co/SkVuien0t8
_PurpleUnicorns|twitter|0.0|0.0|1.0|0.0|RT @l4444k: Snoop Dogg @ Donald Trump Roast https://t.co/SkVuien0t8
NannyDiaries|AbbeWright|0.0|0.0|1.0|0.0|"RT @AbbeWright: When I was canvassing to #GOTVforHRC yesterday, a 4-year-old told me ""Donald Trump shouldn't be allowed to be President."" A"
goawayitsnotme|terrie_ralston|0.0|0.0|1.0|0.0|RT @terrie_ralston: We voted Trump!  #FoxNews2016
MazurekPaul|Pamela_Moore13|-0.4199|0.157|0.843|0.0|"RT @Pamela_Moore13: Trump voter turn-out is way up, polls proven to be rigged. It's happening! https://t.co/6ug1lm0wzZ"
MazurekPaul|twitter|-0.4199|0.157|0.843|0.0|"RT @Pamela_Moore13: Trump voter turn-out is way up, polls proven to be rigged. It's happening! https://t.co/6ug1lm0wzZ"
DrGonzalezH1|ClarkCountyNV|0.0|0.0|1.0|0.0|RT @ClarkCountyNV: Trump campaign petition asks to preserve early voting records. This is required by state law &amp; so it is something we are
mauisrf7|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
mauisrf7|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
shernandez227|themoneygame|0.5719|0.0|0.821|0.179|RT @themoneygame: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/RTr54mdgR3 https://t.co/y
shernandez227|businessinsider|0.5719|0.0|0.821|0.179|RT @themoneygame: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/RTr54mdgR3 https://t.co/y
mallorykrenk|damnnnmoll|0.0|0.0|1.0|0.0|RT @damnnnmoll: I'd rather a cucumber be president instead of trump or hillary
obafan6|LOL_Donkaments|0.0|0.0|1.0|0.0|RT @LOL_Donkaments: #PanHandle GET OUT THERE AND GET #TRUMP IN THE WHITE HOUSE!!!!!!
bulldog338|breitbart|0.6124|0.0|0.75|0.25|Pat Caddell on 'Whatever It Takes': Trump Wins Because 'The People Want Their Country Back' - Breitbart https://t.co/Trn5jjA6P9
HippyMica|40oz_VAN|0.5719|0.0|0.821|0.179|RT @40oz_VAN: How are you leaving the country if Trump wins if you've never even left your city?
karlableal|daanthedevil|0.6597|0.0|0.803|0.197|"RT @daanthedevil: If you vote trump today make sure to explain to your gay, trans, female, Latin, black, and muslim friends why they don't"
jpavlovic801|lottiewillis|-0.4019|0.13|0.87|0.0|"RT @lottiewillis: Insane police presence in Manhattan, right near the Hilton where Trump will be tonight. #ElectionNight #USADecides @newsc"
bbs_firstfed|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
kuyacv|Deadspin|0.0|0.0|1.0|0.0|RT @Deadspin: The Trump campaign wants to make names of Nevada poll workers public. Judge's response: https://t.co/tes99IMbbH
kuyacv|twitter|0.0|0.0|1.0|0.0|RT @Deadspin: The Trump campaign wants to make names of Nevada poll workers public. Judge's response: https://t.co/tes99IMbbH
bisexuaImurphy|sethbeIIamy|0.5423|0.0|0.8|0.2|RT @sethbeIIamy: imagine giving birth to a baby after carrying it for 9 months only for it to become a trump supporter https://t.co/eWAYrhB
bisexuaImurphy|t|0.5423|0.0|0.8|0.2|RT @sethbeIIamy: imagine giving birth to a baby after carrying it for 9 months only for it to become a trump supporter https://t.co/eWAYrhB
DrThomasPaul|DrThomasPaul|0.4199|0.0|0.878|0.122|RT @DrThomasPaul: This #gay woman will tell you like it is. To the #gays brainwashed by #MSM: #WakeUP! #Hillary/#gmo #Trump #LGBTQhttps://
taedybear1230|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
taedybear1230|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
danarose1022|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
heatcost245780|MichaelCBender|-0.3724|0.124|0.876|0.0|RT @MichaelCBender: TRUMP VOTERS:*16% say he's not qualified to serve*18% say he doesn't have effective temperament*13% would be concern
_tylerdurbin|Advil|0.3818|0.0|0.867|0.133|@Advil I would love to keep 90% of America from voting but I'm not part of the Trump campaign.
_ALEXXXXX__|kinkytchalla|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
_ALEXXXXX__|twitter|0.4404|0.0|0.873|0.127|RT @kinkytchalla: Good morning everyone including Eric trump who can go to jail for up to a year for posting this https://t.co/E6WdD70gch
kitsterart|LOLGOP|0.0516|0.138|0.714|0.148|RT @LOLGOP: EXIT POLL: 3 in 10 Trump supporters had trouble finding the exit to the polls.
chased022212|twitter|-0.75|0.444|0.556|0.0|What a freaking idiot. Go trump! #ElectionNight #Election2016 #FoxNews2016 #MakeAmericaGreatAgain https://t.co/Bqn0W6ocRr
ArxipovNifont|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
ArxipovNifont|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
cellydoumerc|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
janakatharine8|hollywoodreporter|0.4019|0.0|0.856|0.144|RT TheRyanParker: These #TrumpCake memes are going to help us all get through the night: https://t.co/ZFm9wlUfNm  https://t.co/AcALMa6TJS
monsungatan|Telegraph|-0.3818|0.115|0.885|0.0|"RT @Telegraph: Now, if somebody cant handle a Twitter account, they cant handle the nuclear codes. Obama Trump losing Twitter access #E"
GetYouAStace|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
GetYouAStace|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
blueefoxxx|mikethenice1|0.0|0.0|1.0|0.0|"RT @mikethenice1: As The Election Comes To A Close, Turnout At Trump Rallies Is Massive https://t.co/wfwytJir8F"
blueefoxxx|westernjournalism|0.0|0.0|1.0|0.0|"RT @mikethenice1: As The Election Comes To A Close, Turnout At Trump Rallies Is Massive https://t.co/wfwytJir8F"
kensiemitchelll|twitter|0.5719|0.0|0.575|0.425|thankful for KY and Trump  https://t.co/zxVvGmpe1i
nousgnostic|PeterSweden7|0.0|0.0|1.0|0.0|"RT @PeterSweden7: So far with votes counted in IN, KY &amp; NH:Trump: 149 808 (68%)Clinton: 62 250 (28%)#ElectionNight"
DaniiT13|HillaryClinton|0.3182|0.0|0.867|0.133|"RT @HillaryClinton: ""Nobody respects women more than me."" Donald TrumpOther things he's said about women: https://t.co/fM9h1WYHkK"
DaniiT13|twitter|0.3182|0.0|0.867|0.133|"RT @HillaryClinton: ""Nobody respects women more than me."" Donald TrumpOther things he's said about women: https://t.co/fM9h1WYHkK"
Jackel_Ramzilla|paulbirkett3|0.3612|0.0|0.894|0.106|RT @paulbirkett3: Choosing between Clinton and Trump to run a nation is like choosing between jimmy saville and the McCanns to babysit your
SpookyHoracio|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
SpookyHoracio|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
rstruglia17|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
rstruglia17|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
RealLifeChino|DonJuancho__|-0.2263|0.168|0.719|0.114|@DonJuancho__ true but no one wants Donald trump to become president. I'd rather Hillary
Kijwii|yvezayntIaurent|-0.5423|0.22|0.78|0.0|"RT @yvezayntIaurent: white person: idk whos worse: hillary or trumplgbtq, women, black people, immigrants, muslims: trump iswhite pers"
brezypoint|BreitbartNews|0.4019|0.0|0.722|0.278|RT @BreitbartNews: Let your yes be yes... https://t.co/IwvjrrpXun
brezypoint|breitbart|0.4019|0.0|0.722|0.278|RT @BreitbartNews: Let your yes be yes... https://t.co/IwvjrrpXun
Civil_war_elect|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: In the two FL counties I've been following, Trump is DRAMATICALLY outperforming Obama from 2012."
sbarrack785|DaRealDanBaulch|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
sbarrack785|t|-0.6705|0.256|0.744|0.0|"RT @DaRealDanBaulch: ""Donald Trump leads by example, closely poll watching as a suspected illegal immigrant attempts to vote."" https://t.co"
jamieraegomes|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
jamieraegomes|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
dovmontagafono2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
dovmontagafono2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
blancbeatz|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: Report: President George W. Bush didn't vote for either Trump, Clinton. #ElectionNight #FoxNews2016 https://t.co/wKkrha8Bqn"
blancbeatz|twitter|0.0|0.0|1.0|0.0|"RT @FoxNews: Report: President George W. Bush didn't vote for either Trump, Clinton. #ElectionNight #FoxNews2016 https://t.co/wKkrha8Bqn"
__naturallylala|chelseahandler|0.3612|0.0|0.906|0.094|"RT @chelseahandler: Stevie Wonder said that voting for Trump is like asking me to drive."" Id rather have Stevie as my Uber driver than Tr"
Smajor1995|AdamYT|0.9195|0.042|0.601|0.357|"@AdamYT @Seapeekay i find it so weird how like all the other states can vote trump, but if hillary gets like CA, NY, FL, WA, OH she wins ha"
DannyChallenger|TrumpBritain|0.0|0.0|1.0|0.0|RT @TrumpBritain: BREAKING NEWS: NEW EXIT POLLTRUMP UP 2% nationally.THE LAND SLIDE IS COMING.RT! RT! Time to #draintheswa
nickwills20|Dan_Siman|0.5719|0.0|0.802|0.198|"RT @Dan_Siman: Let's be real guys, if Trump wins, you are not moving to another country"
GinoVelez201|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
pridbor5|JoePrich|0.1189|0.146|0.693|0.162|RT @JoePrich: Until the polls close in the battlegrounds the media is going to act like Trump is losing baaaaad. So just be prepared
MssLiberty|LyleKlich|-0.4588|0.2|0.8|0.0|RT @LyleKlich: Nevada Poll Workers Break Law: Caught Wearing 'Defeat Trump' T-Shirts https://t.co/ITtwENhUU2
MssLiberty|thegatewaypundit|-0.4588|0.2|0.8|0.0|RT @LyleKlich: Nevada Poll Workers Break Law: Caught Wearing 'Defeat Trump' T-Shirts https://t.co/ITtwENhUU2
TerriMathes|Breaking911|-0.6705|0.256|0.744|0.0|RT @Breaking911: PHOTOS: Trump Tower Surrounded By Dump Trucks Filled With Sand To Edge Against Attacks - TMZ https://t.co/DxcqUSuIXT
TerriMathes|twitter|-0.6705|0.256|0.744|0.0|RT @Breaking911: PHOTOS: Trump Tower Surrounded By Dump Trucks Filled With Sand To Edge Against Attacks - TMZ https://t.co/DxcqUSuIXT
rogdotjpg|Cain_Unable|0.0|0.0|1.0|0.0|"RT @Cain_Unable: I just tried to Vote Trump &amp; the staff wouldn't let me just because I'm ""in Kent"" &amp; ""this is a Tesco self service checkout"
CaseyHill23|twitter|-0.5423|0.538|0.462|0.0|fuck donald trump https://t.co/ZgaROyKXeS
jamie_kerlin|brujaaverde|-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
jamie_kerlin||-0.5859|0.16|0.84|0.0|RT @brujaaverde: Trump couldn't even vote for himself because his mother was born in Scotland you past-ripe banana lookin bitch https://t.c
theriseofgomez|vibeeeez|-0.5574|0.261|0.739|0.0|RT @vibeeeez: prediction: Hillary Clinton is our next present &amp; everyone is shocked Trump lost
actindia|DipDhingani|0.9091|0.0|0.55|0.45|"RT @DipDhingani: #Trump might win the election, but #Modi won the hearts. Haha. #blackmoney #FightAgainstCorruption #OnThisDay #CurrencyB"
Legochanful|GameTheoryRejct|-0.2323|0.193|0.652|0.155|RT @GameTheoryRejct: Meta Theory: Donald Trump will win the election WITH THE POWER OF THE CHAOS EMERALDS?! https://t.co/44jaJJ7Joq
Legochanful|twitter|-0.2323|0.193|0.652|0.155|RT @GameTheoryRejct: Meta Theory: Donald Trump will win the election WITH THE POWER OF THE CHAOS EMERALDS?! https://t.co/44jaJJ7Joq
angel_kat_|u8387p8800|0.0|0.0|1.0|0.0|What a clown. https://t.co/MRKvf1q9Ex
pyrocreativeart|twitter|0.8398|0.0|0.5|0.5|"Let's all pray for Trump, think positive and keep the faith! https://t.co/ESoWNvbGh0"
AlisonLayell|LarrySchweikart|-0.5423|0.2|0.8|0.0|"RT @LarrySchweikart: Trump likely to pick up +40,000 in Brevard alone, 27,000 in Pasco. R counties crushing it, Panhandle already @ 80%R@ 5"
Ceewelsh|BernieSanders|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Ceewelsh|iwillvote|-0.7351|0.396|0.478|0.126|RT @BernieSanders: I hope today we defeat Donald Trump and we defeat him badly. https://t.co/8ttsSwcsnl https://t.co/4Q1JDdglhV
Citizen_USA1|KellyannePolls|0.7096|0.0|0.781|0.219|RT @KellyannePolls: Trump Campaign &amp; RNC @Reince hand in glove. This is about GOP elected officials bragging they voted 3rd party or skippe
misshome888|mitchellvii|0.5719|0.0|0.85|0.15|"RT @mitchellvii: Romney won Brevard County by 36,000 votes in 2012.  I calculate Trump leads it by 52,000 votes.  +16,000 votes for Trump o"
benavi10|WeLoveRobDyrdek|0.4404|0.0|0.791|0.209|RT @WeLoveRobDyrdek: Jon Stewart and Donald Trump beef is funny af https://t.co/j1HsilMOlH
benavi10|twitter|0.4404|0.0|0.791|0.209|RT @WeLoveRobDyrdek: Jon Stewart and Donald Trump beef is funny af https://t.co/j1HsilMOlH
oldschoolvet74|viralnewsx|0.6523|0.1|0.651|0.249|"RT @viralnewsx: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://t.c"
oldschoolvet74||0.6523|0.1|0.651|0.249|"RT @viralnewsx: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://t.c"
bevJacks|SimonNRicketts|0.0|0.0|1.0|0.0|"RT @SimonNRicketts: ""At last, I can finally tweet this. Donald Trump is a  https://t.co/mqk7DWlLSL"
bevJacks|twitter|0.0|0.0|1.0|0.0|"RT @SimonNRicketts: ""At last, I can finally tweet this. Donald Trump is a  https://t.co/mqk7DWlLSL"
teresarc17|michellerj1019|0.0|0.0|1.0|0.0|"RT @michellerj1019: Trump leads Clinton by 120,000 votes  the first Republican candidate to EVER lead in early voting in Florida. #Electio"
angellbadass|BalmainBoslick|-0.1027|0.065|0.935|0.0|RT @BalmainBoslick: Everybody keep askin who I'm voting for idk Hillary gon take my Guns &amp; Trump gon take my FoodStamps
ponyopoundcake|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
rharrisonfries|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana 0.5% reporting TRUMP 70.1% | Hillary 26.1% massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Electi
vivien091011|HaskelBiz|0.5277|0.0|0.714|0.286|"@HaskelBiz @DonaldJTrumpJr I vote Trump, give him a chance. I Can't let her fool me twice "
dionisiyaovchi8|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
dionisiyaovchi8|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
Down4Sue|AdelleNaz|0.0|0.0|1.0|0.0|"RT @AdelleNaz: Star-Spangled Banner being sung by diverse group of Americans in front of #HiltonMidtown, where Trump-Pence ElectionNight pa"
KazakovaAnetta|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
KazakovaAnetta|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
golubev_gektor|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
golubev_gektor|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
jlo4422|FoxNewscomments|0.0|0.0|1.0|0.0|@FoxNewscomments made by KArl Rowe about Trump's comments about G. Bush shouldn't have been allowed-polls haven't closed across the U.S.
NoUghhh|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
HumanMalteser|FrankJavCee|-0.7277|0.63|0.37|0.0|@FrankJavCee Trump!!! FUCK #CrookedHillary
alexisbahl1603|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Liverpotlian|joshgroban|0.6996|0.0|0.799|0.201|"RT @joshgroban: Last night Trump said "" vote tomorrow for all your dreams to come true"" and ""this is our Independence Day!"" He went from Pe"
michaeljohns|pavoterservices|0.0|0.0|1.0|0.0|#Pennsylvania:Polls close at 8pm ET (in one hour). Find your polling location here:https://t.co/5wa27WJ8z1#TrumpPA #TrumpTrain #Trump
ericfrancois19|MadelnCanada|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
ericfrancois19|twitter|0.0|0.0|1.0|0.0|RT @MadelnCanada: #MeanwhileInCanada if Trump wins.. #ElectionNight https://t.co/MzLXBdjcXh
EmilVelour|mitchellvii|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
EmilVelour|t|0.8176|0.0|0.694|0.306|"RT @mitchellvii: In numerous exits, people said they most wanted a change candidate. Trump wins on change 82-12%  Wow. https://t.co/shd8wGO"
harrysuckszayn|TheFunnyVine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
harrysuckszayn|vine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
Donna72Miller|kurteichenwald|0.5984|0.0|0.85|0.15|"RT @kurteichenwald: What I just saw unfold in Nevada with ""Trump v. Hispanics Who Voted"" was some of the most remarkable minutes in a court"
Dre_NoOvO|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
wavvycee|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
wavvycee|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
argiolv|Cam_Major|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
argiolv|twitter|-0.8074|0.477|0.523|0.0|"RT @Cam_Major: ""Trump you a bitch ass nigga and i hope...."" https://t.co/4JDMo5nlWq"
KaitoMelt|twitter|0.5719|0.0|0.575|0.425|USA if #Trump wins. #electionday https://t.co/tNZqUZqFKA
florbarbiebitch|YouTube|0.4753|0.0|0.764|0.236|I liked a @YouTube video from @roiwassabi https://t.co/9WeKnzEHzF DONALD TRUMP IS ILLUMINATI! | Akinator
florbarbiebitch|youtube|0.4753|0.0|0.764|0.236|I liked a @YouTube video from @roiwassabi https://t.co/9WeKnzEHzF DONALD TRUMP IS ILLUMINATI! | Akinator
JimnBL|jaketapper|0.3566|0.0|0.894|0.106|"RT @jaketapper: But then Trump couldn't run, since his mom and paternal grandparents weren't born in the US. So, um, yeah. https://t.co/7Ux"
JimnBL|t|0.3566|0.0|0.894|0.106|"RT @jaketapper: But then Trump couldn't run, since his mom and paternal grandparents weren't born in the US. So, um, yeah. https://t.co/7Ux"
sweetviolets1|HRC4Prison|0.0|0.0|1.0|0.0|"RT @HRC4Prison: Watch out for hoaxes calling Trump's website racist/sexist/etc. Trump website has code flaw, allows you to put whatever h"
hazelstacyyy_|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
zaurav|JYSexton|-0.6874|0.294|0.706|0.0|"RT @JYSexton: If Trump freaks out and destroys the Trump Cake, this whole thing still wasn't worth it but..."
benni_tweets|LordAshcroft|0.0|0.0|1.0|0.0|RT @LordAshcroft: Early US exit polls. Georgia Trump +3. Virginia Clinton+8. N. Carolina Clinton+2. Ohio Tie. Florida Clinton +2. New Hamps
MartinGianolla|VanityFair|0.0772|0.0|0.925|0.075|RT @VanityFair: Even businesses renting space in Trumps landmark building have tangled with the billionaire https://t.co/LbXf329MEX https:
MartinGianolla|vanityfair|0.0772|0.0|0.925|0.075|RT @VanityFair: Even businesses renting space in Trumps landmark building have tangled with the billionaire https://t.co/LbXf329MEX https:
dcutler1958|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
dcutler1958|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
Brainykid2010|twitter|0.7412|0.0|0.786|0.214|"NC, Amer needs your help! This is an elec abt Amer! I appeal to U 2 put country FIRST! Help us to rid our gov of th https://t.co/Ry9CL6cqA3"
Toxlcityy|twitter|0.0|0.0|1.0|0.0|"People on my timeline having meltdowns over Kentucky and Indiana going Trump, get a grip, pick up a book https://t.co/irlqiuFF29"
richardlee_tn|TheRyanParker|0.4019|0.0|0.863|0.137|RT @TheRyanParker: These #TrumpCake memes are going to help us all get through the night: https://t.co/oiuXDIrSf9 #electionday https://t.co
richardlee_tn|hollywoodreporter|0.4019|0.0|0.863|0.137|RT @TheRyanParker: These #TrumpCake memes are going to help us all get through the night: https://t.co/oiuXDIrSf9 #electionday https://t.co
BRIANcates6|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
BRIANcates6|lifezette|0.0|0.0|1.0|0.0|RT @IngrahamAngle: WATCH: @LifeZette is live streaming Donald Trump's remarks now in New York City!Tune in here: https://t.co/6jQdTt7iQm
Giannaamarieeee|owensupertramp|0.2105|0.256|0.407|0.338|RT @owensupertramp: don't mistake my hate for trump with support for hillary. we're either fucked or super weenie hut fucked
vyntage_lo|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
vyntage_lo|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Nicole80017|VictoriaAveyard|0.7269|0.136|0.568|0.297|"RT @VictoriaAveyard: ""It would be sweet sweet justice if it was the Latino vote that stopped Trump."" - Ana Navarro continuing to spit fire."
whitebg19611|TruthAndTime4|0.0|0.0|1.0|0.0|"@TruthAndTime4 you are part of the poorly educated, I see why you are Deplorable! Trump is a Serial Sexual Predator #JustFacts"
spiritofshiloh|"realDonaldTrump,my"|0.0|0.0|1.0|0.0|"#FoxNews2016 I voted 4 @realDonaldTrump,my daughter voted 4 Trump &amp; her doggie Hank is howling for Trump to WIN!Dr https://t.co/bKaR6yzf8D"
spiritofshiloh|twitter|0.0|0.0|1.0|0.0|"#FoxNews2016 I voted 4 @realDonaldTrump,my daughter voted 4 Trump &amp; her doggie Hank is howling for Trump to WIN!Dr https://t.co/bKaR6yzf8D"
brittanynb_|McDanielJustine|0.0|0.0|1.0|0.0|RT @McDanielJustine: Toomey says he voted for trump
bedwcr|ladygaga|0.0|0.0|1.0|0.0|@ladygaga VOTE TRUMP. ONLY REAL PRESIDENT RUNNING THIS ELECTION.
michaelvlueder|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
michaelvlueder|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
Spicedmama|TheView|-0.3089|0.106|0.894|0.0|"RT @TheView: ""I'm a Republican. I don't think Donald Trump is,"" @AnaNavarro says. ""What I see today is not the Republican party . . . that"
queridajesyn|jaw_cee|0.431|0.0|0.898|0.102|RT @jaw_cee: If you're Mexican &amp; voting for Trump let me just say: 1. He doesn't give a fuck about you2. Eres un pendejo3. We don't clai
rivera_chris11|adal_mulero|0.0|0.0|1.0|0.0|@adal_mulero trump arriba
ughxvenus|pettyblackgirI|-0.3612|0.258|0.569|0.174|"RT @pettyblackgirI: After Trump loses tonight, hopefully we'll get more pictures of white ppl crying like they did after Mitt Romney lost t"
rghoover1|realDonaldTrump|-0.25|0.168|0.714|0.117|"RT @realDonaldTrump: 'America must decide between failed policies or fresh perspective, a corrupt system or an outsider'https://t.co/ll8QI"
katepurkis|KathLlewellyn|0.5859|0.0|0.84|0.16|"'even if Trump does win, he has a short attention span so won't be able to concentrate for 4 years in office' @KathLlewellyn"
willddot15|Andy_roodle|0.3612|0.0|0.667|0.333|RT @Andy_roodle: Up like Donald Trump
FreelancerDave|mitchellvii|0.0|0.0|1.0|0.0|RT @mitchellvii: The fact leads are so large in  KY and IN makes me think Trump is getting monster vote and dem crossovers.
RAMSEYUNKNOWN|vox|0.3818|0.0|0.852|0.148|There are 5 people alive who have ever been president. None of them voted for Trump. - https://t.co/AFx6OOLmbR
Bammers05|TBNSport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
Bammers05|tbnsport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
seaexpattrader|reuters|-0.6249|0.24|0.76|0.0|"First U.S. polls close as voters pick between Clinton, Trump after brutal campaign https://t.co/QW5L4qtijD"
TheBreeHive|Cncoll|-0.7003|0.294|0.574|0.132|RT @Cncoll: Not to mention the months of hate speech and fear mongering spewed out by trump. Please be careful tonight.  https://t.co/a1Yur
TheBreeHive|t|-0.7003|0.294|0.574|0.132|RT @Cncoll: Not to mention the months of hate speech and fear mongering spewed out by trump. Please be careful tonight.  https://t.co/a1Yur
lostinthought37|TheFunnyVine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
lostinthought37|vine|0.6369|0.0|0.656|0.344|RT @TheFunnyVine: Still the best Donald Trump vine https://t.co/fPDKVpVnqt
marselmolchano2|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
marselmolchano2|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
RealJoeMirto|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
VEN0MKlNG|GraphicTweetss|-0.6124|0.364|0.636|0.0|RT @GraphicTweetss: Trump = open racistHillary = closet racist https://t.co/6QK3XJe2ID
VEN0MKlNG|twitter|-0.6124|0.364|0.636|0.0|RT @GraphicTweetss: Trump = open racistHillary = closet racist https://t.co/6QK3XJe2ID
Schoroeder|jl095v|-0.5267|0.236|0.764|0.0|RT @jl095v: Can't wait till Obama retard issues gonnneeeeeeeeeeeeeeee go TRUMP  #ElectionNight
YNWAReds96|MenInBlazers|0.3612|0.0|0.839|0.161|RT @MenInBlazers: Trump cake looks like Aaron Ramsey's hair on Arsene Wenger's face https://t.co/BCq3wwmGsM
YNWAReds96|twitter|0.3612|0.0|0.839|0.161|RT @MenInBlazers: Trump cake looks like Aaron Ramsey's hair on Arsene Wenger's face https://t.co/BCq3wwmGsM
Iamnowblue|RalstonReports|0.0|0.0|1.0|0.0|RT @RalstonReports: That was the Trump campaign in a nutshell in that NV court hearing:Unprepared.Loony logic.Lack of knowledge.
MeIAmMomo|TheLifeOfKale|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
MeIAmMomo|t|0.5719|0.0|0.812|0.188|"RT @TheLifeOfKale: Someone said this gone be the national anthem if Trump wins, I'm officially done  https://t.co/MFCsS"
kategoellerr|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
kategoellerr|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
Saeya8|immigrant4trump|0.7506|0.0|0.766|0.234|"RT @immigrant4trump: If you make this go viral, Trump will win. It's about 2 minutes that makes the choice in this election crystal clear h"
Kent_Cyclist|D_Blanchflower|0.0|0.0|1.0|0.0|RT @D_Blanchflower: The name Trump should from this day forward be synonymous with everything we teach our children not to become... 1/2ht
efrosiniyausti7|CrowdFundGurus|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
efrosiniyausti7|reverbnation|0.0|0.0|1.0|0.0|"RT @CrowdFundGurus: Check out ""Donald Trump Your President"" #Trump2016 #TrumpTrain by Rick Poppe - https://t.co/mW0YLUk6aZ"
devery_mccain|twinsational|-0.0258|0.136|0.734|0.13|RT @twinsational: A #Trump Fan Just Pulled A Gun On A Black Voter At #Florida Polling Station - https://t.co/fstiatqr1o
devery_mccain|occupydemocrats|-0.0258|0.136|0.734|0.13|RT @twinsational: A #Trump Fan Just Pulled A Gun On A Black Voter At #Florida Polling Station - https://t.co/fstiatqr1o
globalissuesweb|twib|0.0|0.0|1.0|0.0|America heads to the polls in 2016 elections  as it happened https://t.co/OysLeKsgiF https://t.co/iXgK8Cf0jQ
JEdgar43|ryanjreilly|-0.4588|0.143|0.857|0.0|RT @ryanjreilly: The Trump team says a poll watcher was threatened with a belt. Here's what happened. It's very Philly. https://t.co/c5P3Ex
JEdgar43|t|-0.4588|0.143|0.857|0.0|RT @ryanjreilly: The Trump team says a poll watcher was threatened with a belt. Here's what happened. It's very Philly. https://t.co/c5P3Ex
VGVG0|USATODAY|-0.34|0.13|0.87|0.0|RT @USATODAY: Internet goes crazy over photo of Trump appearing to look at Melania's ballot https://t.co/tmtQvFaeSJ https://t.co/BtkAIIDJFK
VGVG0|usatoday|-0.34|0.13|0.87|0.0|RT @USATODAY: Internet goes crazy over photo of Trump appearing to look at Melania's ballot https://t.co/tmtQvFaeSJ https://t.co/BtkAIIDJFK
