User|Original_User/Web|Compound|Negative|Neutral|Positive|Tweet
HURRICANEPAUL|chelseahandler|0.6369|0.0|0.755|0.245|".@chelseahandler You believed the #FakeNews from @HuffingtonPost that said ""Hillary's chances of winning is 98% to Trump's 2%""LOL#Stupid"
My2cents17|nia4_trump|-0.7184|0.304|0.696|0.0|"RT @nia4_trump: #FridayFeeling Hillary emerged 3 times since her crushing defeat, always wearing purple, the color of Rebellion &amp; Power.  V"
LinBennett|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
GingerJoy98|twitter|0.0|0.0|1.0|0.0|The crazies are running the country. Where are the Dems on Russia hacking?  They need to Benghazi the Republicans l https://t.co/XfzJcpO3aR
tlalmays|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
valfarly|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
BrotherEddy|CNN|-0.4449|0.268|0.732|0.0|@CNN how is Hillary not #1 Hero to CNN?
carolina_brenna|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: What if the election hadn't been hacked?What if Hillary hadn't stole the nomination?What if Obama hadn't given rise to
Llama_Chameleon|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
LVNancy|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
wit_or_whatever|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
smlyc|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
Inked1BNA|Im_ConnorKelley|0.5719|0.0|0.709|0.291|RT @Im_ConnorKelley: @realDonaldTrump @FoxNews Hillary won by 2.83 million votes
jonathanjewel|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
JmyNAMEisJILL|JoelNihlean|0.2263|0.111|0.737|0.152|@JoelNihlean @danfelix82 @justinhendrix @realDonaldTrump This all could have been avoided if Hillary would have been honest about Benghazi.
EpilepticHorse|NotWesleyWelker|-0.296|0.115|0.885|0.0|@NotWesleyWelker @blamemarktjan @PicardTips no the EC is not democratic. T\he people already voted and hillary came out ahead
PatrioticAnnie|Cernovich|0.7717|0.0|0.688|0.312|"RT @Cernovich: Do you trust agents within the CIA, who are Hillary Clinton and Obama loyalists, to tell the truth?"
theidealtwit|asamjulian|-0.5267|0.201|0.738|0.061|"RT @asamjulian: It wasnt Russia, nor Comey. Hillary was an unlikable, uninspiring sociopath w/ no message and multiple legal problems. IT"
nataliedeedah|CronkiteSays|-0.3818|0.205|0.697|0.098|RT @CronkiteSays: REAL NEWSWe've completed an extensive analysis into why Hillary lost and have determined Hillary caused Hillary to lose
DragonPatriota|aqualife2009|0.6597|0.0|0.735|0.265|"@aqualife2009 que se pronuncie Obama SOS malandros. Help us OTAN, help us HillaryAh verdad que gano trump ."
go4gin|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
NorCal_510|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
kingvideo123|RealTimBlack|0.0|0.124|0.714|0.162|"RT @RealTimBlack: Hillary tried to buy the Presidency and failed. Now, how about you tweet about something important like fixing Flint's Wa"
dailydishwater|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
dailydishwater||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
suthernboy100|RepStevenSmith|0.0772|0.0|0.939|0.061|RT @RepStevenSmith: Want to hear about what Hillary did in Libya from a real journalist? @wikileaks Julian Assange explains it in 2 minutes
kcbaseballer50|CarmineZozzora|-0.6705|0.208|0.792|0.0|RT @CarmineZozzora: Fake news narrative check:Russia is to blame for the fact that Hillary and the DNC and the MSM are completely corrupt
badger3030|America_1st_|-0.6901|0.222|0.778|0.0|"RT @America_1st_: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candi"
Fitz5studio|YouTube|0.0|0.0|1.0|0.0|Anonymous   The End Of Hillary Clinton! https://t.co/lofaZIdnMx via @YouTube
Fitz5studio|youtube|0.0|0.0|1.0|0.0|Anonymous   The End Of Hillary Clinton! https://t.co/lofaZIdnMx via @YouTube
laughingat|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
laughingat|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
lowki76|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
lowki76|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
lillyloveyy|patriotrising|-0.4767|0.205|0.795|0.0|The real reason Hillary Clinton is scolding Americans over fake news https://t.co/qlWn81p1Pq https://t.co/stxQbWKtbq
SurvivorMed|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
SurvivorMed|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
clw4packers|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
clw4packers|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
PaschalII|emptywheel|-0.296|0.167|0.833|0.0|"@emptywheel For no reason, today I remembered this piece from primary season  https://t.co/beW9wSxjHG"
PaschalII|pajiba|-0.296|0.167|0.833|0.0|"@emptywheel For no reason, today I remembered this piece from primary season  https://t.co/beW9wSxjHG"
ntvnyr173|naniof_two|0.0|0.0|1.0|0.0|RT @naniof_two: @_edwardmondini_ @ntvnyr173 How about someone start with SOS term + find $6 BILLION Hillary lost/donated to #ClintonFoundat
babysgramma|StevenReyCristo|-0.3425|0.217|0.658|0.124|@StevenReyCristo @Nori_NYCThere is nothing childish about bashing Hillary. She's a liar and a traitor
thereallcherico|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
VozdeRaquel|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
erinpastore|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
Fern0947|reckless_mind|-0.3182|0.095|0.905|0.0|"@reckless_mind @TIME Move to California and bring Hillary with you, then go for walks on trails with her, apparently Secret Service is awol."
Kimmerjo64|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
Kimmerjo64|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
gpnavonod|GodandtheBear|-0.7044|0.272|0.728|0.0|RT @GodandtheBear: What about we don't want Hillary don't you understand? Try all you want you can't make me feel shame for her loss ever.
JIanoale|matthew1nelson1|-0.4019|0.249|0.642|0.109|"@matthew1nelson1 Trump used you. No jobs, no wall, &amp; no jailing Hillary.  He told supporters recently I don't need your votes anymore."
brownlegal|benschwartzy|-0.5177|0.218|0.66|0.122|"RT @benschwartzy: It only took one FBI agent to ruin Nixon (Felt) and one to ruin Hillary (Comey). So, I'm very happy to see Trump making a"
Hay09317403Paul|_News_Trump|-0.6221|0.281|0.719|0.0|RT @_News_Trump: Forget Russia! Reince Priebus Just Pointed Out Why Hillary Really Lost! https://t.co/n8Igft8KNF https://t.co/W2ygPJAJbI
Hay09317403Paul|usapoliticstoday|-0.6221|0.281|0.719|0.0|RT @_News_Trump: Forget Russia! Reince Priebus Just Pointed Out Why Hillary Really Lost! https://t.co/n8Igft8KNF https://t.co/W2ygPJAJbI
c38372346|CarolineWalkerB|-0.4472|0.247|0.629|0.124|"RT @CarolineWalkerB: Hillary Whines About Fake News, So Rush Runs Special 90-Second Montage Just for Her https://t.co/0wgCVLKSQA https://t."
c38372346|conservativefighters|-0.4472|0.247|0.629|0.124|"RT @CarolineWalkerB: Hillary Whines About Fake News, So Rush Runs Special 90-Second Montage Just for Her https://t.co/0wgCVLKSQA https://t."
TCANewsFeed|twitter|-0.6486|0.261|0.739|0.0|RT Roger Stone: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/O5mkAkf9fM #Trump2016
lidia_lidiadim|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
JerseyBoy323|ANOMALY1|0.5719|0.0|0.791|0.209|@ANOMALY1 @chuck270 @KellyannePolls  Hillary surrogate Chris Matthews is brainless-just still tearing @realDonaldTrump-he won #msnbc idiots.
scandallk|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Yankees66y|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
hartfordwolf|Ian56789|-0.4588|0.13|0.87|0.0|RT @Ian56789: Remember when Russian Hackers forced Hillary to wipe her server after being served with a Congressional Sub Poena to preserve
Patrici01435181|gerfingerpoken|0.0|0.0|1.0|0.0|RT @gerfingerpoken: Enabler Hillarys Actions Speak Louder Than Trumps Words - Flopping Aces - https://t.co/zGKDjKzaBM-  https://t.co/Sl1
Patrici01435181|t|0.0|0.0|1.0|0.0|RT @gerfingerpoken: Enabler Hillarys Actions Speak Louder Than Trumps Words - Flopping Aces - https://t.co/zGKDjKzaBM-  https://t.co/Sl1
SusanSt08942260|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
VonnieR57|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
WSCP2|thedailybeast|-0.743|0.296|0.704|0.0|FLASHBACK: Hillarys State Dept Refused to Brand Boko Haram as Terrorists https://t.co/jPCfobm50I #StopHillary #tcot #tlot #TeaParty #PJNet
mswindy12|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
jakezemp|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
gunsrus7|CDCollector23|0.4549|0.0|0.825|0.175|"@CDCollector23 Hillary had way more foreign support than Trump did. Soros, Saudi, Qatar, and others."
Paolalopez1971|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
Paolalopez1971|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
lisajeannemill1|EvelynWhiteGOP|-0.6166|0.237|0.763|0.0|"RT @EvelynWhiteGOP: WATCH  Hillary Calls For CENSORING Conservatives, Her Plan Is SICK https://t.co/5LMuaUi7Sw https://t.co/yrAQudJEOk"
lisajeannemill1|angrypatriotmovement|-0.6166|0.237|0.763|0.0|"RT @EvelynWhiteGOP: WATCH  Hillary Calls For CENSORING Conservatives, Her Plan Is SICK https://t.co/5LMuaUi7Sw https://t.co/yrAQudJEOk"
bikerbd|AndrewWMullins|-0.466|0.138|0.862|0.0|"RT @AndrewWMullins: Wait, whatt?? The Clinton campaign directly tried to get @morningmika pulled from her show for criticizing Hillary? htt"
jakezemp|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
JeffersonObama|6igyak|-0.743|0.27|0.73|0.0|RT @6igyak: Hillary's body double was jealous so it faked being sick just to get back at her.  #BoltonFalseFlagExcuses
allyssar1|twitter|-0.6478|0.218|0.782|0.0|so wasting money on the recount would change the outcome how exactly...now Hillary lost twice and you justify it ho https://t.co/oIXlxFHihM
danieltobin|redsteeze|0.0|0.0|1.0|0.0|RT @redsteeze: Russia wanted Trump. You know who else wanted Trump? Hillary &amp; our media. All three got what they wanted.
wolfy1169|GaetaSusan|-0.8594|0.399|0.498|0.103|"RT @GaetaSusan: Dems, McCain &amp; Graham STOP spreading FAKE NEWS! Every Country hacked Hillary's Private Server! Blame Russia?? What about bl"
Carlene_Meyers|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
Carlene_Meyers|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
rockshout|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
RejectIdolatry|JackPosobiec|-0.7184|0.231|0.769|0.0|"RT @JackPosobiec: Russia didn't cause Hillary to lose the entire Rust Belt and every swing state, her party's failed policies of socialist"
rabiasquared|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
rabiasquared|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
ProgressiveJill|USDefenseWatch|-0.4588|0.267|0.733|0.0|"RT @USDefenseWatch: Hillarys High Drag, Low Speed Campaign Cost a Whopping $1.2Billion https://t.co/Eo8Zi1PqoY https://t.co/J6wjcGfchx"
ProgressiveJill|usdefensewatch|-0.4588|0.267|0.733|0.0|"RT @USDefenseWatch: Hillarys High Drag, Low Speed Campaign Cost a Whopping $1.2Billion https://t.co/Eo8Zi1PqoY https://t.co/J6wjcGfchx"
stickyfacts|mobile|-0.2263|0.213|0.787|0.0|Hillary pleads to dismiss lawsuit against her https://t.co/9ciL3nu3bc
hartzfeld_rick|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Luminami_|realDonaldTrump|-0.7096|0.286|0.656|0.058|@realDonaldTrump Offense is defense. Being offense towards criminal Hillary which still needs her investigation now that they all need to go
d_a_keldsen|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
beckys1girl|MMFlint|-0.6966|0.2|0.8|0.0|RT @MMFlint: Have you heard a ONE Dem leader scream about this? Imagine if Cuba hacked in to throw the election to Hillary? What would Repu
Millenniumistic|brashsculptor1|-0.3318|0.183|0.817|0.0|"RT @brashsculptor1: Seriously, give ONE valid reason Hillary is not now our legal, duly elected PRESIDENT!Welcome, #PresidentClinton "
VonnieR57|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
TheHardMan21|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
wolverines_dad|DailyCaller|-0.5267|0.268|0.614|0.118|RT @DailyCaller: Some Hillary Clinton Donors Infuriated They Didnt Make The Cut For Thank-You Party https://t.co/P7eNNGThpl https://t.co/7
wolverines_dad|dailycaller|-0.5267|0.268|0.614|0.118|RT @DailyCaller: Some Hillary Clinton Donors Infuriated They Didnt Make The Cut For Thank-You Party https://t.co/P7eNNGThpl https://t.co/7
PaxRoHannah|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
jakezemp|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: The Democrats all debate who's going to get out of Hillary's way first, except for VERMONT'S OWN BERNIE SANDERS, who...get"
tparkatheist|directory|0.0|0.0|1.0|0.0|The Atheist in the Trailer Park  : Episode 130: Hillary and the Working Class https://t.co/jAyyOIVicX
inallfandoms|hillyanne23|0.0|0.0|1.0|0.0|RT @hillyanne23: I remember before high school everyone called me Hillary and now all I ever hear is Hill/Hilly and it makes me soooooo hap
whatnext20|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
nanrod98|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
nanrod98||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
exponuntmalum|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
healthygirl90|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
lozanosunwest|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
besthealthever|kr3at|0.0|0.0|1.0|0.0|Michigan Recount: Over 1/2 of Hillary Clintons Detroit Vote Faces Disqualification https://t.co/77DQD6rUhf via @kr3at
besthealthever|alexanderhiggins|0.0|0.0|1.0|0.0|Michigan Recount: Over 1/2 of Hillary Clintons Detroit Vote Faces Disqualification https://t.co/77DQD6rUhf via @kr3at
ConnieBee16|hrtablaze|-0.872|0.405|0.595|0.0|@hrtablaze Hillary lost because she was woefully unsuited for the job. No other reason you pathetic grasping at straws simpletons.
Paolalopez1971|LindaSuhler|0.4404|0.0|0.847|0.153|RT @LindaSuhler: A good time to mention Hillary Clinton's REAL link to Russia...#RussianHackingShe transferred our uranium to Putin...FOR
Millenniumistic|brashsculptor1|-0.5797|0.277|0.61|0.113|RT @brashsculptor1: Nearly 3 million more votes &amp; no cheating. #Hillary is my president.I will accept NOTHING less!#PresidentClinton
Patrici01435181|gerfingerpoken|-0.34|0.179|0.714|0.107|RT @gerfingerpoken: (IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.
Patrici01435181|investors|-0.34|0.179|0.714|0.107|RT @gerfingerpoken: (IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.
Luminami_|realDonaldTrump|-0.1531|0.117|0.789|0.094|"@realDonaldTrump Attack Obama like you did to Hillary Clinton during your speeches. If you say it, it happens. He is moving against you."
Griot_Prince|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
EnigmaNetxx|KatieWagnerFox|0.3818|0.134|0.634|0.231|"RT @KatieWagnerFox: Seth Rich narc'd DNC emails because of cheating in Primary to promote Hillary. #SethRich, ultimate Bernie Bro, RIP. #"
ManyaZuba|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
ManyaZuba|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
GlennOstrosky|realDonaldTrump|-0.6166|0.268|0.732|0.0|RT @realDonaldTrump: HILLARY FAILED ALL OVER THE WORLD. #BigLeagueTruth  LIBYASYRIAIRANIRAQASIA PIVOTRUSSIAN RESETBENGHAZI#D
lks62|terrij68|-0.3317|0.106|0.894|0.0|RT @terrij68: @KellyannePolls almost 3 million more Americans voted for Hillary!!! Most do not want him or at this point you either
westontnicoll|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
AMike4761|America_1st_|-0.6901|0.222|0.778|0.0|"RT @America_1st_: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candi"
mountain_viper|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
nanaz1|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/ynLdIxTaHV
tparkatheist|trailerparkatheist|0.0|0.0|1.0|0.0|Episode 130: Hillary and the Working Class https://t.co/vwNAz6UtJh
RobieCur|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
RobieCur|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
DaFiendR|umpire43|-0.5859|0.137|0.863|0.0|RT @umpire43: Hundreds of thousands of Fraud Hillary votes were foung in Detroit and in Millwaukee and in Philly. Did Russia do that to hel
DanielDastti|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
Cubannator|twitter|0.5859|0.0|0.78|0.22|You mean the Democrats that continue funding tyrants like Castro who beat Cubans daily? Please remind Hillary she l https://t.co/A2cfAkGhi0
jinouyang|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
GigiB84|Harry1T6|0.0772|0.11|0.769|0.121|RT @Harry1T6: Impressive how Russian hackers forced Hillary Clinton to say she would put coal miners out of business and raise their taxes.
TimpoAndante|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
321Chapp|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
321Chapp|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
MicheleWeiss69|mitchellvii|0.0|0.0|1.0|0.0|"@mitchellvii @TRUMP_PREZ what I don't understand...is why the focus isn't on what Hillary did, but how we found out."
Patta47cake|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
zoyeahhhh|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
PatreciaRogers|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
PatreciaRogers|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
RobertTripp12|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
DaVinciVerita|RepStevenSmith|0.0772|0.0|0.939|0.061|RT @RepStevenSmith: Want to hear about what Hillary did in Libya from a real journalist? @wikileaks Julian Assange explains it in 2 minutes
CruzinAhead|SteveDeaceShow|0.0|0.0|1.0|0.0|"RT @SteveDeaceShow: Can only imagine what some ""conservatives"" would say if President Hillary's SOS was a corporate globalist seen toasting"
BitcoinPaul|Freshoutoftissu|0.2716|0.152|0.621|0.227|@Freshoutoftissu @bradmillscan @kazonomics @TheNewBTCGuy @Lunar_Trader no one fucking cares about Hillary.
egopanthers|DonaldsAngel|-0.3182|0.173|0.827|0.0|RT @DonaldsAngel: .@asamjulian .@LindaSuhler .@mitchellvii .@Cernovich .@JackPosobiec Hillary Lost because #ItWasHer@DonaldsAngel https:/
egopanthers||-0.3182|0.173|0.827|0.0|RT @DonaldsAngel: .@asamjulian .@LindaSuhler .@mitchellvii .@Cernovich .@JackPosobiec Hillary Lost because #ItWasHer@DonaldsAngel https:/
Mark_David2|ThePatriot143|-0.4215|0.318|0.682|0.0|@ThePatriot143  he lies as much as hillary
An0nKn0wledge|twitter|-0.5859|0.16|0.84|0.0|They Told Me I Couldn't Have Aliens Hillary &amp; Election Fraud In Same Tweet It Couldn't Be Done They We're Wrong.. https://t.co/ZOOpjH9KmN
Byrlyne|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
boxcoach_dan|baileylewis23|0.0258|0.0|0.95|0.05|@baileylewis23 @stranahan  Assad is  opposed to the pipeline. Investors are the ones trying to oust him. It's why the arabs backed Hillary
Nolanelle|mobile|-0.2263|0.119|0.881|0.0|Hillary pleads court to dismiss lawsuit against her4her lies&amp;harm RE#Benghazi https://t.co/h8Qe9bvVxY. #ImWithHer #StillWithHer #tcot #cvot
Luminami_|realDonaldTrump|-0.4767|0.124|0.876|0.0|@realDonaldTrump Do not be quiet. Speak of the voting machines changing votes from Hillary to Trump. All her votes were yours. Attack them.
JkbComic|twitter|-0.4717|0.128|0.872|0.0|Ken is just another Globalist Hillary Shill who is Butthurt That his Crook HRC didn't Win so that she could carry o https://t.co/Nx8iGaAz5P
Konamali1|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
Konamali1|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
suzost|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
suzost|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
michaelirwin57|Bencjacobs|-0.5688|0.187|0.813|0.0|"@Bencjacobs Based on the history of this current administration, I believe that more then a conspiracy theory the R https://t.co/P9CuN4dCNO"
michaelirwin57|twitter|-0.5688|0.187|0.813|0.0|"@Bencjacobs Based on the history of this current administration, I believe that more then a conspiracy theory the R https://t.co/P9CuN4dCNO"
BongBong|TheRealDonnacha|0.5267|0.0|0.764|0.236|@TheRealDonnacha @bobbyrobertspdx @jowrotethis Right because Hillary was such a fabulous human being: https://t.co/bOjeI7Z9QD
BongBong|youtube|0.5267|0.0|0.764|0.236|@TheRealDonnacha @bobbyrobertspdx @jowrotethis Right because Hillary was such a fabulous human being: https://t.co/bOjeI7Z9QD
gerfingerpoken2|americanthinker|-0.7269|0.357|0.643|0.0|Petraeus Prosecuted - Why not Hillary 4 the same crime? https://t.co/2nLmcsZPVO   - American Thinker - #PJNET - https://t.co/rSFqkggtoF
georgezab|CitizensFedUp|0.2023|0.0|0.872|0.128|"RT @CitizensFedUp: Hillary could have legal right to challenge electoral college system and be next US president, says law professor https:"
paulbenedict7|manny_ottawa|-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
paulbenedict7||-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
lngawaitedsleep|CrankyEthicist|0.7409|0.0|0.773|0.227|"@CrankyEthicist @meakoopa GAME THEORY: MARIO IS ACTUALLY OBAMA, BOWSER IS HILLARY???PARAKOOPA IS THE LOVABLE MEME GUY FROM THE DEBATES"
TheRichWilkins|twitter|-0.6652|0.28|0.72|0.0|"Hillary had an ""email issue"" based on fuzzy conspiracy theories, but the CIA is clueless? https://t.co/h19rVi5ulB"
ericsusy|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
ericsusy|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
DJSCHEMES|twitter|0.0|0.0|1.0|0.0|"""You know I voted for hillary too my nigga"" https://t.co/RK1QDhs4qB"
Markperugini1|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
DonTrumpeone|LindaSuhler|0.4404|0.0|0.847|0.153|RT @LindaSuhler: A good time to mention Hillary Clinton's REAL link to Russia...#RussianHackingShe transferred our uranium to Putin...FOR
john_brumjo|Old_Bern_Kenobi|-0.7579|0.255|0.745|0.0|RT @Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of fac
kmy17|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
DeRay_Shawn|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
CuAtSea|VegasGOP|-0.7778|0.244|0.756|0.0|RT @VegasGOP: Maybe Hillary lost because she is one of the most hated and corrupt individuals to ever seek the Presidency? #AMJoy https://t
CuAtSea||-0.7778|0.244|0.756|0.0|RT @VegasGOP: Maybe Hillary lost because she is one of the most hated and corrupt individuals to ever seek the Presidency? #AMJoy https://t
christiang415|IdiotDems|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
christiang415|t|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
zztopf450|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
zprfct|phil200269|-0.875|0.348|0.576|0.076|RT @phil200269: Hillary getting on the fake news bandwagon is like Bill Clinton speaking out against the evils of rape in American society.
1stworldmusic|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
ShockedBirgit|BV|0.0|0.0|1.0|0.0|The misjudgments about voters began with Hillary Clinton's announcement video. https://t.co/29SvDZiVeA via @BV #StillSanders
ShockedBirgit|bloomberg|0.0|0.0|1.0|0.0|The misjudgments about voters began with Hillary Clinton's announcement video. https://t.co/29SvDZiVeA via @BV #StillSanders
Trippn21|jojoh888|-0.5574|0.419|0.581|0.0|@jojoh888 And #Hillary shit her pants
leelamchop|DailyCaller|-0.5267|0.268|0.614|0.118|RT @DailyCaller: Some Hillary Clinton Donors Infuriated They Didnt Make The Cut For Thank-You Party https://t.co/P7eNNGThpl https://t.co/7
leelamchop|dailycaller|-0.5267|0.268|0.614|0.118|RT @DailyCaller: Some Hillary Clinton Donors Infuriated They Didnt Make The Cut For Thank-You Party https://t.co/P7eNNGThpl https://t.co/7
filmystic|zachheltzel|0.3182|0.079|0.722|0.199|"RT @zachheltzel: 68% of Trump supporters want him to imprison Hillary Clinton for no reason, in case you were wondering the exact number of"
thiaalife|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
lrnewton1|RNRMississippi|-0.2263|0.215|0.642|0.143|"RT @RNRMississippi: Russians are Amazing: Set up a private server, rigged the primary, used BleachBit to violate a court order, then made"
naniof_two|_edwardmondini_|0.0|0.0|1.0|0.0|@_edwardmondini_ @ntvnyr173 How about someone start with SOS term + find $6 BILLION Hillary lost/donated to #ClintonFoundation!
ReGenesisRadio|youtube|0.3724|0.045|0.852|0.103|https://t.co/shE8LxIjnF it's not the Russians stupid its the NSA and FBI Hillary they don't want you in there get a clue zip go away u2 BHO
alohaberni|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
hillary_sarah|tatianaramozzzz|0.0|0.0|1.0|0.0|@tatianaramozzzz kkkkkkkk Jesus
TXhistorylover|twitter|-0.25|0.125|0.875|0.0|The Russians replicated every voter in America and cancelled all of the Hillary votes https://t.co/RC7GpYkJyR
mauriciod44|riwired|0.2023|0.0|0.921|0.079|"RT @riwired: Pres. Obama sent his top campaign manager, and other aides, on American taxpayer $ to influence Israel's election &amp; Hillary in"
extractionista|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
test5f1798|nydailynews|0.0|0.0|1.0|0.0|https://t.co/yv4h9sR6iN : f4b96ade-2c88-4500-b802-11c64292b1ad
CerulloElaine|bfraser747|-0.6901|0.222|0.778|0.0|"RT @bfraser747:  ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."" ~ @GovMikeHu"
suzierwilson|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
gretchen_nation|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
aasstevens|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
kgiuseppe|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/FRzp92uwwv via @Change
kgiuseppe|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/FRzp92uwwv via @Change
SukiFrench|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
PatriciaAHenso1|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
MLinebacker48|MarieLeff|-0.4767|0.262|0.611|0.127|RT @MarieLeff: @BreitbartNews This is better than the daily reminder that Hillary suffered a brain injury so severe... 
MrDevilAdvocate|RNRMississippi|-0.2263|0.215|0.642|0.143|"RT @RNRMississippi: Russians are Amazing: Set up a private server, rigged the primary, used BleachBit to violate a court order, then made"
hillary_sarah|tatianaramozzzz|0.0|0.0|1.0|0.0|RT @tatianaramozzzz: @hillary_sarah serissimo kkjkkkkkkk
kgvet|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
jjwright_janet|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
go4gin|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
tatianaramozzzz|hillary_sarah|0.0|0.0|1.0|0.0|@hillary_sarah serissimo kkjkkkkkkk
Barbara4Freedom|SteveDeaceShow|0.0|0.0|1.0|0.0|"RT @SteveDeaceShow: Can only imagine what some ""conservatives"" would say if President Hillary's SOS was a corporate globalist seen toasting"
02C5|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
PeteKaliner|redsteeze|0.0|0.0|1.0|0.0|RT @redsteeze: Russia wanted Trump. You know who else wanted Trump? Hillary &amp; our media. All three got what they wanted.
MarkopoloXYZ|davidfrum|0.0|0.0|1.0|0.0|"RT @davidfrum: Maybe it wasnt tactical, but I still dont understand why Hillary never said: Take off that pin, its not your flag, you P"
grocknroll165|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
HaieyEHampton|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
techweenie|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
yceek|yceek|0.0|0.0|1.0|0.0|"RT @yceek: Americans! If Hillary Clinton can stage assassin of Trump in Reno, imagine what this thug do to the rest of us! https://t.co/Ed"
yceek|t|0.0|0.0|1.0|0.0|"RT @yceek: Americans! If Hillary Clinton can stage assassin of Trump in Reno, imagine what this thug do to the rest of us! https://t.co/Ed"
Dupetones|camper_bruce|0.0|0.0|1.0|0.0|@camper_bruce @thehill Hillary slept thru Hillary's part
wilmajeanne|morningmika|-0.5423|0.29|0.71|0.0|@morningmika @JoeNBC @MSNBC @HillaryClinton @chucktodd @jasoninthehouse You warned us Hillary.  Unfortunately e-mai https://t.co/TZAvJtWY2T
wilmajeanne|twitter|-0.5423|0.29|0.71|0.0|@morningmika @JoeNBC @MSNBC @HillaryClinton @chucktodd @jasoninthehouse You warned us Hillary.  Unfortunately e-mai https://t.co/TZAvJtWY2T
Beatromney|AdamsFlaFan|-0.3612|0.167|0.739|0.094|"RT @AdamsFlaFan: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/wokIcX3tph via @crooksandliars"
Beatromney|crooksandliars|-0.3612|0.167|0.739|0.094|"RT @AdamsFlaFan: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/wokIcX3tph via @crooksandliars"
imalilr|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
texan2you|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
texan2you|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
1AllHearingEar|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
Inked1BNA|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
GGthinking|slone|-0.4466|0.118|0.882|0.0|RT @slone: We KNOW that McCain and Graham voted for Hillary b/c they're both GLOBALISTS. There is NO difference btwn a D globalist &amp; an R g
vandives|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
michellegun24|umpire43|-0.5859|0.137|0.863|0.0|RT @umpire43: Hundreds of thousands of Fraud Hillary votes were foung in Detroit and in Millwaukee and in Philly. Did Russia do that to hel
noturbone|hrh_orchid|-0.6808|0.219|0.781|0.0|@hrh_orchid @ybbkaren derp she still lost 30 out of 50 states that means more than 50% of the states rejected hillary clinton
NotTurnbull|peterdaou|-0.25|0.152|0.738|0.111|"RT @peterdaou: If you're convinced that Hillary is corrupt, flawed, unlikable, dishonest, that was EXACTLY the goal of Russian tampering. C"
valfarly|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
ericsusy|DineshDSouza|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
ericsusy|twitter|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
GregQ42|SethAMandel|0.0|0.0|1.0|0.0|"You know what, Democrats?#Hillary cost Hillary the election. Get over it@SethAMandel @seanmdav"
Yombe|theatlantic|-0.5267|0.207|0.793|0.0|The Danger of Trump and Putin's Relationship - The Atlantic9/21/16 #TrumpPutin #Russianhackers #Hillary #Mandate https://t.co/08FyWaCoxI
GoldAntiquated|NIRPUmbrella|0.2942|0.0|0.905|0.095|RT @NIRPUmbrella: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http
stormyzcrochet|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/HYANNDPcxe
mom2kidz63|DineshDSouza|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
mom2kidz63|twitter|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
Therealrajeshp|steph93065|-0.5455|0.144|0.799|0.057|@steph93065 I think they are getting Hillary for 2020 (it's not hillarys fault but Russia) vote for her in 2020 and oh there was fake news.
njpcnjpc|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
GADiA_tx|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
CzarCache_|twitter|0.0|0.0|1.0|0.0|o#dank #memes #meme #fazeup  #fazeclan #crazy #funny #hillary #trump #rattpack #lol #omg #clown #clowns #youtube https://t.co/LVJcs5uD0d
Anyshka|MrDane1982|0.1007|0.161|0.714|0.125|"RT @MrDane1982: 40 yrs of fighting for us, this time we fight for her until she have enough ground to stand on! The best thing Hillary can"
JimmyForTrump|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
YaBoyKentucky|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
YaBoyKentucky|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
masonkiana3|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
masonkiana3|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
chirprn|AdamParkhomenko|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
chirprn|nydailynews|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
torrHL|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
national_newsb|truthfeed|-0.5319|0.186|0.814|0.0|This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/xzYcgnSEdh #RETWEEETME https://t.co/yZ4qa8HVNO
jstacks248|GopAaron|0.5574|0.0|0.566|0.434|@GopAaron thank god crooked Hillary didn't get elected .
shellyhawthorne|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
valfarly|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
VelvaDStevenson|BourneInTexas|-0.34|0.138|0.862|0.0|"RT @BourneInTexas: Tony Blair, Hillary Clinton, Kuwait....and the secret transfer of fundsbut let's blame Russia instead.@Nigel_Farag"
veggie64_leslie|SinCityCarol|-0.4767|0.22|0.78|0.0|RT @SinCityCarol: @veggie64_leslie @HuffPostPol oh for fucks sake. #1 is Hillary herself
DeltaBravoNews|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
DeltaBravoNews|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
jkatsalis|dandrezner|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
jkatsalis|t|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
leezalotte|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
masayanmk2|TrinityNYC|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
masayanmk2|t|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
LisaCBlair|twitter|-0.5562|0.473|0.527|0.0|Put Hillary in prison!   https://t.co/l8bNt6scJe
DagnyDelinquent|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
DagnyDelinquent|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
Lonestar2003|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
RanaeMayle|larryelder|-0.4215|0.258|0.595|0.147|"RT @larryelder: There's no point in a California recount. Hillary won by over 5 million dead people, I mean votes.#Recount2016 https://t."
RanaeMayle||-0.4215|0.258|0.595|0.147|"RT @larryelder: There's no point in a California recount. Hillary won by over 5 million dead people, I mean votes.#Recount2016 https://t."
Jwalkertide|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
Mexicanpov|Mexicanpov|0.0656|0.167|0.658|0.175|"RT @Mexicanpov: LOL, there is So Much wrong doing there, however, in 90mins of pleading his case to DJT in exchange for no pardon of hillar"
lidia_lidiadim|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
lidia_lidiadim|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
kidaisinyou|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
ElisaPerezG1|Ian56789|-0.4588|0.13|0.87|0.0|RT @Ian56789: Remember when Russian Hackers forced Hillary to wipe her server after being served with a Congressional Sub Poena to preserve
RandallBeard88|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
Shawna_08|trumpwallnow|0.0|0.0|1.0|0.0|RT @trumpwallnow: I just found what I'm getting Hillary for Christmas. They come in different colors to match her jumpsuits!https://t.co/v
Shawna_08|abhinavvadrevu|0.0|0.0|1.0|0.0|RT @trumpwallnow: I just found what I'm getting Hillary for Christmas. They come in different colors to match her jumpsuits!https://t.co/v
MissMindfield|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
ThomasT72388202|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
extractionista|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
extractionista|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
ICANFLA|BizPacReview|-0.4019|0.119|0.881|0.0|"Dem gov. of Virginia recalls omen that spelled doom for Hillary, and it has to do with his https://t.co/WjrPjy4qfw  via @BizPacReview"
ICANFLA|bizpacreview|-0.4019|0.119|0.881|0.0|"Dem gov. of Virginia recalls omen that spelled doom for Hillary, and it has to do with his https://t.co/WjrPjy4qfw  via @BizPacReview"
valfarly|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: The Democrats all debate who's going to get out of Hillary's way first, except for VERMONT'S OWN BERNIE SANDERS, who...get"
blueskymountain|DenbrotS|0.25|0.105|0.74|0.155|RT @DenbrotS: IS TRUMP'S DEAL WITH PUTIN THE BIGGEST PAY TO PLAY OF ALL TIME?@realDonaldTrump @oreillyfactor https://t.co/VlNBARG9CS
blueskymountain|linkis|0.25|0.105|0.74|0.155|RT @DenbrotS: IS TRUMP'S DEAL WITH PUTIN THE BIGGEST PAY TO PLAY OF ALL TIME?@realDonaldTrump @oreillyfactor https://t.co/VlNBARG9CS
LCSCHOPP|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
LCSCHOPP|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
jataylor11|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
windwens|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
graydaygamer|lhfang|-0.6908|0.251|0.749|0.0|RT @lhfang: This guy works for David Brock as a partisan pro-Hillary media critic. And just makes shit up. https://t.co/l3LVbndNDK
graydaygamer|twitter|-0.6908|0.251|0.749|0.0|RT @lhfang: This guy works for David Brock as a partisan pro-Hillary media critic. And just makes shit up. https://t.co/l3LVbndNDK
2kschumacher|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
vhhcjhv|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
SSNjl|RepStevenSmith|0.0772|0.0|0.939|0.061|RT @RepStevenSmith: Want to hear about what Hillary did in Libya from a real journalist? @wikileaks Julian Assange explains it in 2 minutes
NewEnglandDevil|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
f77a9c24c7f9451|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
roqchrisy|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
Razorback40|lillyslolly|0.6369|0.0|0.851|0.149|@lillyslolly I watch it all both sides. That's why I can't stand trump or Hillary. But you love to lump everyone into one group or the other
emilypassey|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
ericserati68|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
ericserati68|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
hypnocoach183|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
GmaPeace2|twitter|0.6597|0.0|0.787|0.213|Amazed it's ok with you foreign power commited espionage to put Trump in. If it was Hillary they helped? You'd be s https://t.co/ywnIAaPk1g
EdenVision|gatses13|-0.4278|0.193|0.706|0.101|RT @gatses13: Rush Limbaugh Plays Montage Of Hillary As A Purveyor Of FAKE NEWS https://t.co/JFAGeK9L5I via @YouTube
EdenVision|youtube|-0.4278|0.193|0.706|0.101|RT @gatses13: Rush Limbaugh Plays Montage Of Hillary As A Purveyor Of FAKE NEWS https://t.co/JFAGeK9L5I via @YouTube
realtonydetroit|GeorgeTakei|-0.7783|0.342|0.658|0.0|@GeorgeTakei You are another mindless liberal that is a walking contradiction. Hillary received MILLIONS from Russia. Where's your criticism
02C5|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
jondoepolitics|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
jondoepolitics|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
aallaart|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
ConorOGinger|benschwartzy|-0.5177|0.218|0.66|0.122|"RT @benschwartzy: It only took one FBI agent to ruin Nixon (Felt) and one to ruin Hillary (Comey). So, I'm very happy to see Trump making a"
jonburtonhx|manny_ottawa|-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
jonburtonhx||-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
DanaSlechta66|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
Wayne5Juan|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
SuccessAtEnron|jharlen00|-0.3976|0.309|0.691|0.0|@jharlen00 @vandercyrus @CNN so you blame Hillary
RamBoPirate|HispanicsTrump|0.0|0.0|1.0|0.0|RT @HispanicsTrump: If Hillary really wants to know who cost her the election all she needs to do is look in the mirror... #FakeNews #Russi
mariaso1200|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
MackNDaly|WaukeshaGOP|0.9437|0.055|0.41|0.535|"@WaukeshaGOP I am in no way a hillary supporter, but had to laugh at your spelling... hiLlar? Haha xD"
JamieAgathaRose|twitter|0.0516|0.0|0.845|0.155|"You backed Hillary, you backed these people. Why should we listen to you? https://t.co/4zEHMP82PE"
elizabethkap|BuzzFeedNews|-0.4767|0.181|0.819|0.0|"RT @BuzzFeedNews: Hillary Clinton Calls On Congress, Silicon Valley To Address Fake News Epidemichttps://t.co/poWhi5ZMMY https://t.co/Vy"
elizabethkap|t|-0.4767|0.181|0.819|0.0|"RT @BuzzFeedNews: Hillary Clinton Calls On Congress, Silicon Valley To Address Fake News Epidemichttps://t.co/poWhi5ZMMY https://t.co/Vy"
twodog711|EylinHurt|-0.4824|0.164|0.836|0.0|"RT @EylinHurt: FBI ASST. DIRECTOR COMES OUT, Says HILLARY SHOULD BE SHOT BY FIRING SQUAD https://t.co/HqfWHjakOr https://t.co/bm5Hk5uLbc"
twodog711|conservativefighters|-0.4824|0.164|0.836|0.0|"RT @EylinHurt: FBI ASST. DIRECTOR COMES OUT, Says HILLARY SHOULD BE SHOT BY FIRING SQUAD https://t.co/HqfWHjakOr https://t.co/bm5Hk5uLbc"
stiNgo100|theGSpledge|-0.3889|0.26|0.601|0.139|@theGSpledge @kestans NO you lie. Hillary did not PBO did not. Your anger is hurting you.
JohnBlast2000|johncitysq|-0.2023|0.162|0.714|0.124|"RT @johncitysq: Do you, @elliottkrista, remember Dems said anyone concerned over election integrity was a ""Threat to Democracy""?https://t."
JohnBlast2000||-0.2023|0.162|0.714|0.124|"RT @johncitysq: Do you, @elliottkrista, remember Dems said anyone concerned over election integrity was a ""Threat to Democracy""?https://t."
carterdsc|gerfingerpoken2|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
carterdsc|americanthinker|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
geno2u|realDonaldTrump|-0.128|0.131|0.757|0.112|@realDonaldTrump @NBCNightlyNews @CNN Were they trashing Hillary again. Sick of hearing she is way ahead by millions in the popular vote.
emilypassey|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
emilypassey||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
michellegun24|RNRMississippi|-0.2263|0.215|0.642|0.143|"RT @RNRMississippi: Russians are Amazing: Set up a private server, rigged the primary, used BleachBit to violate a court order, then made"
Stupidosaur|Stupidosaur|-0.802|0.265|0.735|0.0|"RT @Stupidosaur: GST &amp; Aadhaar are part of same scam to destroy India's economy, federalism, welfare and democracy. The 'magic wand' Hillar"
macbeezy411|KD_Marshall|0.34|0.0|0.833|0.167|@KD_Marshall @TulsaPolice im assuming you voted for hillary..well you lost..congrats you played yourself
SenSlomkowski|twitter|-0.2411|0.197|0.803|0.0|Didn't you endorse Hillary Clinton? Now that's hypocrisy. https://t.co/JhHEAYMBJg
TlyaShontal|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
dunnkath|terrij68|-0.3317|0.106|0.894|0.0|RT @terrij68: @KellyannePolls almost 3 million more Americans voted for Hillary!!! Most do not want him or at this point you either
jcschmieder|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
FisherBurton|BillyVonElds|0.0|0.0|1.0|0.0|@BillyVonElds Address my tweets about Hillary first. You haven't yet.
jumba47|kurteichenwald|-0.2382|0.22|0.67|0.11|"RT @kurteichenwald: No offense, @chucktodd, but when u say no one was sure Russia behind hack pre-election, shows u need to read more. http"
DTParallelogram|hillary_square|0.0|0.0|1.0|0.0|@hillary_square @RhombusGary @KiteBernie @JillRectangle @TrapezoidTed I know that quads should have opposite sides that are congruent
Azrosco|tteegar|-0.3182|0.095|0.905|0.0|RT @tteegar: .@PrisonPlanet Libtards b likeHow many ways can we rub a historic Hillary Clinton loss in &amp; pour salt on this wound we con
JamesS020770|AmericanMex067|-0.6486|0.22|0.735|0.045|"RT @AmericanMex067: She had fake news backing her, DOJ, Obama - spent $1.2 billion &amp; still lost. Russia had nothing 2 do w/it.https://t.co"
Miitomoan|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
LiliaMorraz|ThreatcoreNews|-0.4019|0.213|0.787|0.0|RT @ThreatcoreNews: .@smerconish I guess the Russians hacked Hillary's crowds too? #investigate
Ranthruredlight|MtnMD|0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
Ranthruredlight||0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
euriag|TecReview|0.0|0.0|1.0|0.0|RT @TecReview: As fue como Donald Trump pudo superar a Hillary Clinton en los ltimos das de campaa en Estados Unidos https://t.co/7dgPZ
euriag|t|0.0|0.0|1.0|0.0|RT @TecReview: As fue como Donald Trump pudo superar a Hillary Clinton en los ltimos das de campaa en Estados Unidos https://t.co/7dgPZ
mowser1970|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
di8285502|DaveH_RPh|0.0|0.0|1.0|0.0|@DaveH_RPh are those the Hillary voters?
ntvnyr173|_edwardmondini_|0.0|0.0|1.0|0.0|RT @_edwardmondini_: @ntvnyr173   Hillary would be a female version of Carter.......on steroids.
pauIrevere|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Pallamus|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
Pallamus|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
GigiB84|amrightnow|0.0|0.0|1.0|0.0|RT @amrightnow: Hillary Clinton should be in Jail Not on the campaign Trail #realdonaldtrump #military #army #navy #usmc https://t.co/6VIfN
GigiB84|t|0.0|0.0|1.0|0.0|RT @amrightnow: Hillary Clinton should be in Jail Not on the campaign Trail #realdonaldtrump #military #army #navy #usmc https://t.co/6VIfN
crossfitnans|crossfitnans|0.0|0.0|1.0|0.0|RT @crossfitnans: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/dEI2GxZF5y via @Change
crossfitnans|change|0.0|0.0|1.0|0.0|RT @crossfitnans: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/dEI2GxZF5y via @Change
PerryBullock|redsteeze|0.0|0.0|1.0|0.0|RT @redsteeze: Russia wanted Trump. You know who else wanted Trump? Hillary &amp; our media. All three got what they wanted.
allofusfortrump|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
dierdremccormic|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
dierdremccormic|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
RiseUpAbove|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
kgvet|BarrieNJ|0.6322|0.0|0.794|0.206|RT @BarrieNJ: The Nate Silver that predicted Hillary would win in a monumental landslide?  That Nate Silver? https://t.co/nUaXgBN3aB
kgvet|twitter|0.6322|0.0|0.794|0.206|RT @BarrieNJ: The Nate Silver that predicted Hillary would win in a monumental landslide?  That Nate Silver? https://t.co/nUaXgBN3aB
AnxietyMisfit|OddLane|0.0|0.0|1.0|0.0|RT @OddLane: The First Amendment as suggestion box: https://t.co/jQ45zepGyP #HillaryClinton #Fakenews
AnxietyMisfit|reason|0.0|0.0|1.0|0.0|RT @OddLane: The First Amendment as suggestion box: https://t.co/jQ45zepGyP #HillaryClinton #Fakenews
mtduarte_|MadameWoo69|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
mtduarte_|change|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
emilypassey|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
djjohnso|emptywheel|0.0|0.0|1.0|0.0|@emptywheel @majorajam this article from UPI was a week or two after Conway took over. She understood this effect https://t.co/TrCL7CIDop
djjohnso|upi|0.0|0.0|1.0|0.0|@emptywheel @majorajam this article from UPI was a week or two after Conway took over. She understood this effect https://t.co/TrCL7CIDop
PxlJedi|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
bd05926|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
thecatsmeow0410|Old_Bern_Kenobi|-0.7579|0.255|0.745|0.0|RT @Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of fac
JackieGlo305|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
3Panda3|NotJoshEarnest|0.0|0.0|1.0|0.0|RT @NotJoshEarnest: Hillary tried to go to Wisconsin and Michigan but the Russians kept hacking her plane back to California and New York
Trumps1stMember|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
Pab1oFresh|SouthPark|-0.5267|0.139|0.861|0.0|"these @SouthPark trump/hillary episodes not only show how f*ed up their politics are, it shows how f* stupid the writers are #boycott"
1ofabev|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
suzykq5|KailiJoy|0.0|0.0|1.0|0.0|"RT @KailiJoy: Anyway. You can expect that I'll be talking about Hillary Clinton, the president who should have been, for the next four year"
wooofpak987|igob4u2|-0.2481|0.117|0.817|0.066|"RT @igob4u2: #ECvoteHRC 12/19 @HillaryClinton Have you signed #ElectoralCollegePetition? Plz do! Need 6 mil signs, Stuck at 4.8 https://t.c"
wooofpak987||-0.2481|0.117|0.817|0.066|"RT @igob4u2: #ECvoteHRC 12/19 @HillaryClinton Have you signed #ElectoralCollegePetition? Plz do! Need 6 mil signs, Stuck at 4.8 https://t.c"
mikew6161|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
Michael01466880|farathomas|0.0|0.0|1.0|0.0|"@farathomas @steph93065 the Democrats fixing the primaries,media tilting polls towards Hillary, crooked media  investigate that"
national_newsb|thefederalistpapers|-0.3182|0.173|0.827|0.0|Why R#ussia Had NOTHING To Do With Hillarys Loss https://t.co/C2eYqXBeFV #RETWEEETME https://t.co/Lij8NiW8ga
qtelektra|FrankLuntz|-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
qtelektra||-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
GoodwinHH6|dachsiemoron|0.0|0.0|1.0|0.0|RT @dachsiemoron: What did he say about Hillary's? https://t.co/8uHktYC1fx
GoodwinHH6|twitter|0.0|0.0|1.0|0.0|RT @dachsiemoron: What did he say about Hillary's? https://t.co/8uHktYC1fx
GlennOstrosky|realDonaldTrump|-0.5439|0.164|0.836|0.0|RT @realDonaldTrump: Hillary said she was under sniper fire (while surrounded by USSS.) Turned out to be a total lie. She is not fit to lea
AnnTruwe|ArianeBellamar|0.0|0.0|1.0|0.0|RT @ArianeBellamar:  b4 Partisan! Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/CMOS
AnnTruwe|t|0.0|0.0|1.0|0.0|RT @ArianeBellamar:  b4 Partisan! Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/CMOS
Karabee3|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
Karabee3||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
MethodVine|bestofhomer|-0.4767|0.437|0.563|0.0|@bestofhomer hillary knows even worse
burksclaudine1|burksclaudine1|0.5719|0.0|0.764|0.236|RT @burksclaudine1: @WhiteHouse our rights to have a president voted by the people.Hillary won
Politics_Info|politicsinformer|-0.7269|0.379|0.621|0.0|Madonna and Hillary: Witch and Nasty Woman as Sisters inArms https://t.co/qsFHztvwsb https://t.co/gIRIc9noyc
suzykq5|KailiJoy|-0.6007|0.176|0.824|0.0|"RT @KailiJoy: And now Hillary, who gave us everything of herself and never got a thank you, gets to go on all the goddamned makeup-free hik"
Michelem1998|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
COBYKOEHL|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
WriterRx|TheFreeWorld1|-0.4939|0.158|0.842|0.0|RT @TheFreeWorld1: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #WorldHunger https://t.co
WriterRx|t|-0.4939|0.158|0.842|0.0|RT @TheFreeWorld1: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #WorldHunger https://t.co
Cindy63306167|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
Cindy63306167|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
trump1supporter|KellyannePolls|0.0338|0.152|0.626|0.222|"@KellyannePolls @ErengwaM @Newsweek If he did, thank you Putin because Hillary sure as hell didn't go without help as in $1.2 billion spent"
Maritza03239786|NIRPUmbrella|0.2942|0.0|0.905|0.095|RT @NIRPUmbrella: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http
bikerbd|michelekirkBPR|-0.7269|0.336|0.664|0.0|RT @michelekirkBPR: One man in Hillarys campaign warned she could lose and everybody ignored him https://t.co/A1z3VKU2OE https://t.co/Ahda
bikerbd|bizpacreview|-0.7269|0.336|0.664|0.0|RT @michelekirkBPR: One man in Hillarys campaign warned she could lose and everybody ignored him https://t.co/A1z3VKU2OE https://t.co/Ahda
GregQ42|SethAMandel|-0.296|0.115|0.885|0.0|"RT @SethAMandel: ""Russia cost Hillary the presidency"" is another way of saying ""no one I know voted for Trump."""
ginaboyer|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
tonic516|stylistkavin|-0.7269|0.289|0.711|0.0|RT @stylistkavin: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/pqjurgsNw7 #SistersinArms @Madonna @Hillar
tonic516|nytimes|-0.7269|0.289|0.711|0.0|RT @stylistkavin: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/pqjurgsNw7 #SistersinArms @Madonna @Hillar
forte2x|NormOrnstein|-0.395|0.25|0.75|0.0|@NormOrnstein but haven't they promised to continue investigating Hillary?
CattHarmony|redsteeze|0.0|0.0|1.0|0.0|RT @redsteeze: Russia wanted Trump. You know who else wanted Trump? Hillary &amp; our media. All three got what they wanted.
hillary_sarah|tatianaramozzzz|0.0|0.0|1.0|0.0|@tatianaramozzzz srio? 
ntvnyr173|_edwardmondini_|0.0|0.0|1.0|0.0|"RT @_edwardmondini_: @ntvnyr173   Everyone thinks Hillary has all this ""experience"":  would we call Benghazi, Libya, Syria &amp; Russia ""experi"
relevantspur|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
reneeepona|WLTaskForce|-0.4898|0.143|0.857|0.0|@WLTaskForce @christymatson64 @wikileaks @CBSNews Hillary -people with souls see that U sold yours to evil-U lost bc of who you are!!!
Byrlyne|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
TechnicalGuryou|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
TechnicalGuryou|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
crossfitnans|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/dEI2GxZF5y via @Change
crossfitnans|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/dEI2GxZF5y via @Change
lindsayrda53|MelindaThinker|0.2023|0.0|0.833|0.167|RT @MelindaThinker: Russian interference with the election could give courts legal authority to install Hillary https://t.co/By58AeeOe3
lindsayrda53|huffingtonpost|0.2023|0.0|0.833|0.167|RT @MelindaThinker: Russian interference with the election could give courts legal authority to install Hillary https://t.co/By58AeeOe3
ErnstKoby|OttomanZealot|0.0|0.0|1.0|0.0|RT @OttomanZealot: I don't believe Russia was behind the email hacks but you all do realize that those emails were HER emails regardless. H
JoanSebastian__|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
JoanSebastian__|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
Rosamelchoto69|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
Rosamelchoto69|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
Pepitopatea777|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
Pepitopatea777|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
laprofe63|MMFlint|-0.6966|0.2|0.8|0.0|RT @MMFlint: Have you heard a ONE Dem leader scream about this? Imagine if Cuba hacked in to throw the election to Hillary? What would Repu
Phaedrus08|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: Think bout this: Allied intel servives investigating prez-elect 2 learn if he's Putin stooge in place 2 shatter NATO ht
DuckGuyy42|NozNewz_com|-0.5319|0.186|0.814|0.0|RT @NozNewz_com: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/OSGmSmxWoO
DuckGuyy42|linkis|-0.5319|0.186|0.814|0.0|RT @NozNewz_com: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/OSGmSmxWoO
dj4k4000|slone|-0.4466|0.118|0.882|0.0|RT @slone: We KNOW that McCain and Graham voted for Hillary b/c they're both GLOBALISTS. There is NO difference btwn a D globalist &amp; an R g
2figures2|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
2figures2|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
Vote_American|KellyannePolls|0.4389|0.116|0.657|0.228|"@KellyannePolls @DavidWeingust Hillary &amp; Her Entourage are Clearly Out Classed, Outdated &amp; Rude! Maybe U can find them a Safe Place, Jail?"
DTWhitehouseDT|CLIFFBELL888|-0.6486|0.238|0.676|0.085|@CLIFFBELL888 congress defunding security is to blame. likely the same story for the hundreds of dead embassy workers before hillary was SoS
jdraina|JackBPR|-0.6486|0.325|0.675|0.0|@JackBPR @SNL continues to campaign for Hillary. Mocks Trump. Change the channel. Morons.
TheMrsDarcy|syqau|-0.6351|0.224|0.776|0.0|"RT @syqau: During recount, in 100 precincts in Milwaukee, WI,  Hillary Clinton lost 17,000 votes!! (Trump lost only 1,700) https://t.co/VS"
TheMrsDarcy|t|-0.6351|0.224|0.776|0.0|"RT @syqau: During recount, in 100 precincts in Milwaukee, WI,  Hillary Clinton lost 17,000 votes!! (Trump lost only 1,700) https://t.co/VS"
twodog711|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
cckeefe|Mediaite|0.0|0.0|1.0|0.0|RT @Mediaite: Former U.S. Ambassador to Russia: Vladimir Putin Wanted 'Revenge' on Hillary Clinton https://t.co/e4Kfd6FfcB (VIDEO) https://
cckeefe|mediaite|0.0|0.0|1.0|0.0|RT @Mediaite: Former U.S. Ambassador to Russia: Vladimir Putin Wanted 'Revenge' on Hillary Clinton https://t.co/e4Kfd6FfcB (VIDEO) https://
mama2fluffs|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
mama2fluffs|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
jesskivlehen|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
psmccusker|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: #PodestaEmails more proof of Hillary's Russian Connections. ""Grassley Letter"" to Loretta Lynch. #CorruptMedia let this stor"
RickySi16087724|WEdwarda|-0.9466|0.49|0.51|0.0|"RT @WEdwarda: RUSH Limbaugh DESTROYS Hillary With Montage Of LIES In VIRAL VIDEO After She Blamed ""Fake News"" For Her Loss https://t.co/0rm"
RickySi16087724|t|-0.9466|0.49|0.51|0.0|"RT @WEdwarda: RUSH Limbaugh DESTROYS Hillary With Montage Of LIES In VIRAL VIDEO After She Blamed ""Fake News"" For Her Loss https://t.co/0rm"
_edwardmondini_|ntvnyr173|0.0|0.0|1.0|0.0|@ntvnyr173   Hillary would be a female version of Carter.......on steroids.
NLTCNY|Portosj81J|0.2263|0.0|0.924|0.076|RT @Portosj81J: If the CIA knew that Russia was behind hacking then why did Obama allow Hillary to use a private server with official secre
lorilpeabody|HispanicsTrump|0.0|0.0|1.0|0.0|RT @HispanicsTrump: If Hillary really wants to know who cost her the election all she needs to do is look in the mirror... #FakeNews #Russi
Evilmititis|Krisp_y|-0.0059|0.192|0.583|0.225|"RT @Krisp_y: Hillary supporters, as highly hypocritical as you are, please repeat after me: ""Russia didn't rig it, she just lost"" https://t"
Evilmititis||-0.0059|0.192|0.583|0.225|"RT @Krisp_y: Hillary supporters, as highly hypocritical as you are, please repeat after me: ""Russia didn't rig it, she just lost"" https://t"
fransis48|StopStopHillary|0.4019|0.0|0.863|0.137|"RT @StopStopHillary: #Pizzagate's looking real enough to hire a special prosecutor to look into #Weiner, #Podesta, &amp; #Hillary. #SecretCIA h"
WolfNW|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
WolfNW||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
deborahjlundy|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
adjunctprofessr|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
Compact987|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
Compact987|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
g_rubylee2009|MtnMD|0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
g_rubylee2009||0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
InEgo_|twitter|-0.0094|0.229|0.544|0.227|Sure. Obama torpedoed Hillary so that Trump won so that he can blame the Russians and declare war. https://t.co/eoMC1g9Dwm
Eyes_of_justice|USDefenseWatch|-0.4588|0.267|0.733|0.0|"RT @USDefenseWatch: Hillarys High Drag, Low Speed Campaign Cost a Whopping $1.2Billion https://t.co/Eo8Zi1PqoY https://t.co/J6wjcGfchx"
Eyes_of_justice|usdefensewatch|-0.4588|0.267|0.733|0.0|"RT @USDefenseWatch: Hillarys High Drag, Low Speed Campaign Cost a Whopping $1.2Billion https://t.co/Eo8Zi1PqoY https://t.co/J6wjcGfchx"
l_RW_Offen5iveT|twitter|-0.6124|0.273|0.727|0.0|"Egotistical Hillary demanded customized BB when SoS. NSA said no, so she &amp; staff entered SCIFs w insecured devices https://t.co/ICRgIqiLQG"
claramanoucheka|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
claramanoucheka|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
Balthier28|_CillaW|0.2732|0.0|0.92|0.08|RT @_CillaW: Agreed. It's all deep rooted sexism. Imagine if Hillary was elected &amp; doing half of the things Trump is right now. People woul
gregjamesbarton|dandrezner|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
gregjamesbarton|t|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
US_Threepers|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Riley4Reason|jus1_kimberely|-0.6124|0.263|0.737|0.0|@jus1_kimberely @MikeMil84124709 @JudicialWatch @irs None of your accusations against Hillary make Crooked Trump's problems go away.
DA4Liberty|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
149049c1e543418|RepStevenSmith|0.0772|0.0|0.939|0.061|RT @RepStevenSmith: Want to hear about what Hillary did in Libya from a real journalist? @wikileaks Julian Assange explains it in 2 minutes
test5f1798|nydailynews|0.0|0.0|1.0|0.0|https://t.co/yv4h9sR6iN : a03ca8f5-dbc6-4f1b-afb9-64124588998b
kaseymend|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/n3G83XEpMd via @Change
kaseymend|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/n3G83XEpMd via @Change
CeeStarrr|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
digitalorality|socalmike_SD|0.0|0.0|1.0|0.0|RT @socalmike_SD: Wikileaks: Hillary Clinton Bragged About Being Invited to Putin's 'Inner Sanctum' https://t.co/UyYrkL9WlO via @BreitbartN
digitalorality|breitbart|0.0|0.0|1.0|0.0|RT @socalmike_SD: Wikileaks: Hillary Clinton Bragged About Being Invited to Putin's 'Inner Sanctum' https://t.co/UyYrkL9WlO via @BreitbartN
DaleF3|eztempo|-0.6249|0.212|0.788|0.0|@eztempo @CNN I blame Hillary and her DWS campaign manager installed at the DNC. They planned this coronation since her 2008 lose.
Tokaise|johncitysq|-0.2023|0.162|0.714|0.124|"RT @johncitysq: Do you, @elliottkrista, remember Dems said anyone concerned over election integrity was a ""Threat to Democracy""?https://t."
Tokaise||-0.2023|0.162|0.714|0.124|"RT @johncitysq: Do you, @elliottkrista, remember Dems said anyone concerned over election integrity was a ""Threat to Democracy""?https://t."
dms1013|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
Hillarizer|hillaryclinton|-0.0352|0.182|0.645|0.174|"#HillaryWhines About Fake News, So Rush Runs Special 90-Second #MontageJust for Her https://t.co/3o37eH4nXi"
VelvaDStevenson|Tis4Ta|-0.1779|0.182|0.657|0.161|"RT @Tis4Ta: Still no lead in Seth Rich death, he work for the government. They should be looking with a fine tooth comb, But for Hillary ev"
SinCityCarol|veggie64_leslie|-0.4767|0.256|0.744|0.0|@veggie64_leslie @HuffPostPol oh for fucks sake. #1 is Hillary herself
Katja_Thieme|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
SGT_B_Dub|sean_spoonts|0.0|0.0|1.0|0.0|RT @sean_spoonts: This is why Hillary shouldn't have had that private server. All this goes back to that. https://t.co/HniijJKggx
SGT_B_Dub|twitter|0.0|0.0|1.0|0.0|RT @sean_spoonts: This is why Hillary shouldn't have had that private server. All this goes back to that. https://t.co/HniijJKggx
mserna95|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/Sw9nNqT02t via @Change
mserna95|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/Sw9nNqT02t via @Change
rosendo_joe|MaxBlumenthal|0.0|0.0|1.0|0.0|RT @MaxBlumenthal: .@AliAbunimah @JoyAnnReid What we've learned here is that Putin took out Hillary but Hillary did not take out Qaddafi. h
Aszneth|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
Aszneth|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
notrelluf|vivelafra|-0.5251|0.195|0.805|0.0|"@vivelafra @chucktodd He's a MSM lickspittle, but if you think he's a Hillary shill you're fucking nuts."
LivingOn18|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
fk_eduardo|thomaswikjr|0.4019|0.0|0.847|0.153|"@thomaswikjr @Graham1Sam @GodandtheBear Yes. There were two choices, the apocalypse or Hillary. You chose the apocalypse."
MMaria03146111|DCClothesline|-0.7351|0.323|0.677|0.0|RT @DCClothesline: Hillary Clinton  The Queen of Fake News  Lectures Americans About Fake News https://t.co/AlPAn3K3Xc
MMaria03146111|dcclothesline|-0.7351|0.323|0.677|0.0|RT @DCClothesline: Hillary Clinton  The Queen of Fake News  Lectures Americans About Fake News https://t.co/AlPAn3K3Xc
txconservgirl|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
THEscottywilly|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
THEscottywilly|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
election16news|dcexaminer|0.0|0.0|1.0|0.0|@dcexaminer Hillary is in denial. She fell short. #hubris https://t.co/ZJYYNU2fec
election16news|twitter|0.0|0.0|1.0|0.0|@dcexaminer Hillary is in denial. She fell short. #hubris https://t.co/ZJYYNU2fec
Yamil_Sued|regisgiles|-0.2808|0.196|0.666|0.138|QUEEN OF FAKE NEWS: 8 Times Hillary Fabricated Stories to Help Her Image https://t.co/Dx3bWD3n98 via @regisgiles
Yamil_Sued|girlsjustwannahaveguns|-0.2808|0.196|0.666|0.138|QUEEN OF FAKE NEWS: 8 Times Hillary Fabricated Stories to Help Her Image https://t.co/Dx3bWD3n98 via @regisgiles
1carpediem2016|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
allofusfortrump|SenSanders|0.0|0.0|1.0|0.0|@SenSanders  you sold yourself.  You don't count anymore  go back to your Hillary house
MissEMT37|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
s_chelf|idawhannadoyou|-0.1027|0.185|0.69|0.125|RT @idawhannadoyou: (2) hacked #Hillary's mouth forcing her call half of #Trump's supporters deplorable which obviously affected the outcom
thomasfrank1101|reasonedvoices|-0.2732|0.333|0.427|0.239|@reasonedvoices Hillary was asking for war lol
saminhim|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
saminhim|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
SscottSsmith84|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
1baldeagle77|YouTube|0.2732|0.132|0.683|0.185|"Mark Cuban EAT YOUR WORDS, ""Hillary will win the election"", Trump Will Lose https://t.co/rXgMZpCs58 via @YouTube"
1baldeagle77|youtube|0.2732|0.132|0.683|0.185|"Mark Cuban EAT YOUR WORDS, ""Hillary will win the election"", Trump Will Lose https://t.co/rXgMZpCs58 via @YouTube"
thomas_quinlan|catoletters|0.4019|0.0|0.876|0.124|"RT @catoletters: More proof Russians helped Trump.  Russians paid actors to openly support Hillary, knowing that heavily increasd votes for"
scott_stalker2|TerriGreenUSA|-0.0423|0.095|0.818|0.088|"RT @TerriGreenUSA: We've already said no to #fakenews. DSW didn't deny anything wiki said, and there's still the investigation into Hillary"
DirtPacino|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
Volunteerguys|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
SiberiaCat3|cherilyneagar|0.0|0.0|1.0|0.0|.@cherilyneagar MorriseyWV @UrlingTreasurer Hillary: $30B plan to retrain coal workers.  #MoralElectors https://t.co/1xEVHu81gV
SiberiaCat3|huffingtonpost|0.0|0.0|1.0|0.0|.@cherilyneagar MorriseyWV @UrlingTreasurer Hillary: $30B plan to retrain coal workers.  #MoralElectors https://t.co/1xEVHu81gV
Col_Connaughton|youtube|0.0|0.0|1.0|0.0|Hillary Clinton 'FAINTS' At 9/11 Ceremony || RAW FOOTAGE https://t.co/gUVmQettFp #hillary #clinton #faints
NAlejandra2|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Zelidasquare|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
bigdaddydoggie|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
ThorneColleen|nia4_trump|-0.7184|0.304|0.696|0.0|"RT @nia4_trump: #FridayFeeling Hillary emerged 3 times since her crushing defeat, always wearing purple, the color of Rebellion &amp; Power.  V"
psbaloans4u|twitter|0.0|0.0|1.0|0.0|Why would they donate so much money to Hillary lets see how much they donate in 2017 this is plain &amp; simple a https://t.co/zQCQx3R09n
macmc101|CronkiteSays|-0.3818|0.205|0.697|0.098|RT @CronkiteSays: REAL NEWSWe've completed an extensive analysis into why Hillary lost and have determined Hillary caused Hillary to lose
katherinejnowak|teeg_dougland|0.1027|0.0|0.92|0.08|58. pretending sanders didn't contribute to hillary's healthcare attempt as first lady despite obvs proof @teeg_dougland @neeratanden
PolitixGal|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
CBatBG|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
psmccusker|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: Hillary's secret $2.35M Russian Connection was so crooked, even the #CorruptMedia had to covered it. #UraniumOnehttps://t."
lindagknowlton|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
cala_1111|truthfeed|-0.5255|0.195|0.805|0.0|"VIDEO : Rush Limbaugh's New ""Hillary Fake News"" Hit Piece is BLOWING UP the Internet! https://t.co/9hcspkikD1"
NancyPoehler|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
NancyPoehler|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
MaeroCarol|ReaganCoalition|0.0|0.0|1.0|0.0|RT @ReaganCoalition: REVEALED  The Hillary Aide Who KNEW It Was All Over https://t.co/pBxUGkdoYl
MaeroCarol|fiscalconservatives|0.0|0.0|1.0|0.0|RT @ReaganCoalition: REVEALED  The Hillary Aide Who KNEW It Was All Over https://t.co/pBxUGkdoYl
LOPlato|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
CHOCLABLOVER|KailiJoy|-0.872|0.356|0.603|0.041|"RT @KailiJoy: But we want to be lied to. Obviously. And for all the fake scandals and baseless accusations, that's not what Hillary Clinton"
pyalgia|theGSpledge|0.0|0.0|1.0|0.0|"RT @theGSpledge: If there's 1 thing Hillary's disappearance in the face of Trump shows is that she never was a leader, just a self-entitled"
claramanoucheka|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
DDale13|DDale13|-0.5574|0.167|0.833|0.0|@DDale13 Hillary had 22 Ls for the 22 state primaries/caucuses she lost. Clinton has 30 for the 30 states she lost in the general election
MelikaleKamalei|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
LifeisGreat_45|369news|-0.4404|0.195|0.805|0.0|U.N. Official 'Accidentally' Crushes Own Throat Right Before Testifying Against Hillary Clinton https://t.co/EjjoWVO0SI
esparhawk|DineshDSouza|-0.7579|0.365|0.539|0.095|RT @DineshDSouza: .@HillarysAmerica revealed the truth about Hillary and helped avert disaster. Commemorate her historic defeat: https://t.
esparhawk||-0.7579|0.365|0.539|0.095|RT @DineshDSouza: .@HillarysAmerica revealed the truth about Hillary and helped avert disaster. Commemorate her historic defeat: https://t.
bloodinbritish3|GaetaSusan|-0.8594|0.399|0.498|0.103|"RT @GaetaSusan: Dems, McCain &amp; Graham STOP spreading FAKE NEWS! Every Country hacked Hillary's Private Server! Blame Russia?? What about bl"
K_DUBB_80|holistic_pickle|0.7506|0.0|0.769|0.231|"@holistic_pickle ME TOO, TRUMP IS NOT A CONSERVATIVE AT ALL BUT HILLARY TALKED ABOUT HIM NOT RESPECTING THE RESULTS... WELP "
teambernie27001|lhfang|0.743|0.0|0.7|0.3|RT @lhfang: Hillary Clinton as Sec of State created a special division within the agency to promote fracking abroad w/Exxon https://t.co/pA
teambernie27001|t|0.743|0.0|0.7|0.3|RT @lhfang: Hillary Clinton as Sec of State created a special division within the agency to promote fracking abroad w/Exxon https://t.co/pA
SiberiaCat3|stanggt|0.0|0.0|1.0|0.0|.@stanggt @ronestesks Hillary was right again. Dont vote Trump be #MoralElectors https://t.co/P9v6KRqb90 https://t.co/K9f3BUotfD
SiberiaCat3|theguardian|0.0|0.0|1.0|0.0|.@stanggt @ronestesks Hillary was right again. Dont vote Trump be #MoralElectors https://t.co/P9v6KRqb90 https://t.co/K9f3BUotfD
ErengwaM|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
matt_r29|twitter|0.0|0.0|1.0|0.0|#Killary #Hillary has aligned herself as the biggest #LOSER in American history! The people have spoke! https://t.co/nXvCZQljbA
klgillum|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
kellogh|k_villav|-0.284|0.142|0.858|0.0|@k_villav @lpolgreen @chrislhayes it's not a great news source but the Guardian also confirms https://t.co/7R9xdw6unx
kellogh|theguardian|-0.284|0.142|0.858|0.0|@k_villav @lpolgreen @chrislhayes it's not a great news source but the Guardian also confirms https://t.co/7R9xdw6unx
rugratfarm|igob4u2|-0.2481|0.117|0.817|0.066|"RT @igob4u2: #ECvoteHRC 12/19 @HillaryClinton Have you signed #ElectoralCollegePetition? Plz do! Need 6 mil signs, Stuck at 4.8 https://t.c"
rugratfarm||-0.2481|0.117|0.817|0.066|"RT @igob4u2: #ECvoteHRC 12/19 @HillaryClinton Have you signed #ElectoralCollegePetition? Plz do! Need 6 mil signs, Stuck at 4.8 https://t.c"
Kimmerjo64|MADE__USA|-0.6956|0.192|0.808|0.0|RT @MADE__USA: Obama &amp; Hillary where nothing but Political Pickpockets willing to Poison an Entire Country for Billions of Dollars. #Obama
RebelHeartWorld|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
emalone|dandrezner|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
emalone|t|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
reillyzona|MissMandi00|0.0|0.0|1.0|0.0|@MissMandi00 @redcat0827 @peterdaou @tom_kelo And Hillary had a ton of bucks from other foreign powers to counteract that flood.
FishPar4N2|andersonDrLJA|0.5904|0.0|0.832|0.168|RT @andersonDrLJA: I NEVER VOTED 4 #OBAMA; DIDNT VOTE 4 #HILLARY &amp; NEVER WILL; WILL ALWAYS #FIGHTTerrorism; IM PROUD 2B A PATRIOT &amp; FOREVE
riatheo36|ANTI_ALP|0.4048|0.193|0.472|0.335|@ANTI_ALP Hillary is making Rudd look like the world's most gracious loser
LEISUREGODDESS|LeoKapakosNY|-0.6249|0.203|0.797|0.0|RT @LeoKapakosNY: I wonder if @Reince Priebus would have disputed the fact that foreign agents hacked us if it got Hillary elected? I think
johnhashissay|larryelder|-0.4215|0.258|0.595|0.147|"RT @larryelder: There's no point in a California recount. Hillary won by over 5 million dead people, I mean votes.#Recount2016 https://t."
johnhashissay||-0.4215|0.258|0.595|0.147|"RT @larryelder: There's no point in a California recount. Hillary won by over 5 million dead people, I mean votes.#Recount2016 https://t."
khubb64|thehill|-0.4019|0.114|0.886|0.0|@thehill Dems knew Hillary was gonna lose so they set the narrative that someone else caused it. Barack and Hillary caused it.
OurRevolution2|twitter|-0.4939|0.158|0.842|0.0|RT Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failur https://t.co/NWzLrHTaAw
smillr|sean_spoonts|0.0|0.0|1.0|0.0|RT @sean_spoonts: This is why Hillary shouldn't have had that private server. All this goes back to that. https://t.co/HniijJKggx
smillr|twitter|0.0|0.0|1.0|0.0|RT @sean_spoonts: This is why Hillary shouldn't have had that private server. All this goes back to that. https://t.co/HniijJKggx
Huntclub2001|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
Huntclub2001|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
AmericanMom2|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
1sfleming302|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
saucissonsec|joshtpm|-0.4404|0.209|0.791|0.0|@joshtpm @TPM Buuuuuuut... it happened before he was elected and discredited Hillary.
healthygirl90|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
BonnieLCollins3|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
lmpauls51|twitter|-0.4898|0.166|0.834|0.0|"The NSA is ALSO a ""whistleblower"" to keep Hillary OUT of WH! CIA is CNN! Misinformation News! https://t.co/zTfzbn2QAN"
bigdaddydoggie|CelesDavis2|0.4939|0.0|0.868|0.132|@CelesDavis2 @Tablavi @keksalamander @MightyChin Putin has been laughing at Obama &amp; Hillary for 8 years. That is why he does what he wants.
SeminolePost|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
SeminolePost|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
PVan1016|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
alfredanchor|birdistheherd|-0.6124|0.3|0.6|0.1|"@birdistheherd @260a105fb5c7455 Really don't need any lines of attack. Like Hillary, Trump's adversaries usually shoot themself in the foot"
LibrarianTr|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
MuffinAndElliot|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
Dbiggs1007Donna|stopsorosnow|0.5229|0.1|0.718|0.182|@stopsorosnow NO WONDER HILLARY &amp; BILL CLINTON ARE SO TIGHT WITH SOROS! SHE WORSHIPPED SAUL ALINSKY! LOOK AT THE SIMILARITIES BETWEEN THE 2!
healthygirl90|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
Stever0020|Tymeeks98|0.4019|0.0|0.863|0.137|"RT @Tymeeks98: @mitchellvii @JohnFromCranber Didn't Mexico try to help Hillary, by having Mexican citizens infiltrate US election process?"
mikea71|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
hillaryslead|realdonaldtrump.|0.25|0.096|0.735|0.169|"Hillary got 2,841,862 more votes than @realdonaldtrump. Sorry, it's the truth. #nomandate."
NickKruel14|twitter|0.4632|0.101|0.672|0.228|If only Russia didn't hack Hillary's illegal server and leak incriminating emails about her  Seems a lot like Hil https://t.co/UsfWQLumew
EAlfaroQ|billmaher|0.3134|0.048|0.855|0.097|"RT @billmaher: Seeing Hillary speaking yesterday: Thank you, and Bill, for over 30 yrs of service. And now I never want to see either one o"
carpejor512|GeorgeTakei|0.3182|0.0|0.85|0.15|@GeorgeTakei we found out that Hillary supported the fondling of little kids. Much worse.........
Judyjcprov47|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
antonia_nemka|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
WWZ_TAK|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
national_newsb|usapoliticstoday|-0.6221|0.316|0.684|0.0|Forget Russia! Reince Priebus Just Pointed Out Why Hillary Really Lost! https://t.co/4qOJOC21cq https://t.co/hykf8584mN
MyPupVoted|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
SnakePlisskn|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
inradiator|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
MonicaDoss|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
EastOrlandoPost|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
EastOrlandoPost|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
PatPatojson|oguzhan_ciltas|-0.5319|0.177|0.823|0.0|RT @oguzhan_ciltas: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/FbU1BAyxtu https://t.co/67thQUmlZ1
PatPatojson|truthfeed|-0.5319|0.177|0.823|0.0|RT @oguzhan_ciltas: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/FbU1BAyxtu https://t.co/67thQUmlZ1
carolebobarrel|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
nuiotwo|nuiotwo|-0.296|0.241|0.602|0.158|"RT @nuiotwo: Neera Tanden On TPP: ""This Makes Hillary Seem Politically Craven At Best Or A Liar At Worse""  https://t.co/ITyoGUinlI"
nuiotwo|zerohedge|-0.296|0.241|0.602|0.158|"RT @nuiotwo: Neera Tanden On TPP: ""This Makes Hillary Seem Politically Craven At Best Or A Liar At Worse""  https://t.co/ITyoGUinlI"
freewillfighter|gerfingerpoken2|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
freewillfighter|americanthinker|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
LibertySeeds|"LindseyGrahamSC,"|0.34|0.0|0.854|0.146|"#ISIS allies of @LindseyGrahamSC, @Evan_McMullin, and #Hillary #Clinton make gains around #Palmyra, #Syria ... https://t.co/uO4MRdEBU7"
LibertySeeds|zerohedge|0.34|0.0|0.854|0.146|"#ISIS allies of @LindseyGrahamSC, @Evan_McMullin, and #Hillary #Clinton make gains around #Palmyra, #Syria ... https://t.co/uO4MRdEBU7"
healthygirl90|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: The Democrats all debate who's going to get out of Hillary's way first, except for VERMONT'S OWN BERNIE SANDERS, who...get"
JDiviv|youtube|0.0|0.0|1.0|0.0|Putin discusses actions of Obama &amp; HillaryA MUST SEE video:https://t.co/zePLFaDlUa https://t.co/pVGLH1Q2FM
RightAsRain7|rb87700|-0.2732|0.209|0.642|0.15|RT @rb87700: @wolfgangfaustX @WDFx2EU26 @POTUS @Judgenap we were saved from Hillary/DNC/Rino/lying media war w Russia
OrangeTint|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
OrangeTint|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
DorH84607784|realjunsonchan|0.4076|0.133|0.632|0.235|"RT @realjunsonchan: -@KellyannePolls completely rekts Rotten Hillary. Lol. This is how America should be governed, spend less, win more. Ni"
JamesTokarz|YouTube|0.4753|0.0|0.819|0.181|I liked a @YouTube video from @markdice https://t.co/QMRHklItwV Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!
JamesTokarz|youtube|0.4753|0.0|0.819|0.181|I liked a @YouTube video from @markdice https://t.co/QMRHklItwV Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!
saminhim|BarrieNJ|0.6322|0.0|0.794|0.206|RT @BarrieNJ: The Nate Silver that predicted Hillary would win in a monumental landslide?  That Nate Silver? https://t.co/nUaXgBN3aB
saminhim|twitter|0.6322|0.0|0.794|0.206|RT @BarrieNJ: The Nate Silver that predicted Hillary would win in a monumental landslide?  That Nate Silver? https://t.co/nUaXgBN3aB
jlizza1|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
MtnMD|asJBdorightthng|0.0|0.0|1.0|0.0|RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.co/mQwwx3cuBj
MtnMD|occupydemocrats|0.0|0.0|1.0|0.0|RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.co/mQwwx3cuBj
SizzlerKistler|jillybobww|0.3612|0.0|0.912|0.088|RT @jillybobww: It is starting to seem like maybe Hillary's email is the one thing the Russians didn't hack &amp; so we should in fact be askin
amrightnow|twitter|0.0|0.0|1.0|0.0|Hillary Clinton should be in Jail Not on the campaign Trail #realdonaldtrump #military #army #navy #usmc https://t.co/6VIfNZoMGg
Wethepeople196|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: People weren't concerned about Russia when Hillary was selling them US uranium.#MAGA
NorrisImages|gerfingerpoken2|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
NorrisImages|americanthinker|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
1jelliott1|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
MichaelWeschler|mobile|-0.2732|0.204|0.667|0.13|"When you cheat in any race, you're disqualified &amp; the next person wins. Oh, &amp; Hillary has 2.8M more votes. https://t.co/gJ6yPtCwbn #ReVote"
SscottSsmith84|DiamondandSilk|0.0|0.0|1.0|0.0|@DiamondandSilk Bikers For Hillary https://t.co/TripKzLuj0
SscottSsmith84|twitter|0.0|0.0|1.0|0.0|@DiamondandSilk Bikers For Hillary https://t.co/TripKzLuj0
Ariadne38|breitbart|-0.7906|0.438|0.563|0.0|Hillary Clinton: All Rape Victims Deserve To Be Believed - Breitbart https://t.co/WRrDZQrmxe
GeoffDPeterson|dandrezner|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
GeoffDPeterson|t|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
DustyFae|youtube|0.5473|0.0|0.786|0.214|"WANTING ANOTHER ELECTION, HILLARY WILL BE LUCKY TO GET ANY VOTES NEXT TIME https://t.co/gGMP4i7skI"
allyssar1|twitter|0.4374|0.124|0.595|0.28|olo lol I did it I admit it this s why Hillary lost twice llolo boom!! https://t.co/vLoWrJ7uHs
s_chelf|Portosj81J|0.2263|0.0|0.924|0.076|RT @Portosj81J: If the CIA knew that Russia was behind hacking then why did Obama allow Hillary to use a private server with official secre
AuntChellie26|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
Edmundite1|KLSouth|0.0|0.0|1.0|0.0|RT @KLSouth: #ImWithHer #Hillary is yesterday. #FakeNews #SheLost https://t.co/GTIDfrD3in
Edmundite1|twitter|0.0|0.0|1.0|0.0|RT @KLSouth: #ImWithHer #Hillary is yesterday. #FakeNews #SheLost https://t.co/GTIDfrD3in
Mark_David2|Harry1T6|0.0772|0.11|0.769|0.121|RT @Harry1T6: Impressive how Russian hackers forced Hillary Clinton to say she would put coal miners out of business and raise their taxes.
JaynAlexndr|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
bbeekk321|ChipBrooks17|-0.3182|0.113|0.887|0.0|RT @ChipBrooks17: Fact: You can simultaneously believe Hillary lost because America didn't trust/like her while still viewing the Russian h
nightingalern|mobile|-0.3885|0.273|0.727|0.0|HILLARY PLEADS TO DISMISS LAWSUIT AGAINST HER https://t.co/wOm3VZizZ4
ZKondos|INTJutsu|0.5574|0.0|0.833|0.167|@INTJutsu @PatVPeters Merkel did to Germany exactly what Hillary was about to do to the US Thank you God for protecting us the last minute
lugnut4|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
kaiaka|NorthFalcon74|-0.4019|0.114|0.886|0.0|RT @NorthFalcon74: @Portosj81J @Dewblue1 Notice nobody is saying *what* was hacked. The fact is it was Hillary Clinton's server. End of sto
TraceySRogers1|NozNewz_com|-0.5319|0.186|0.814|0.0|RT @NozNewz_com: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/OSGmSmxWoO
TraceySRogers1|linkis|-0.5319|0.186|0.814|0.0|RT @NozNewz_com: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/OSGmSmxWoO
SolUru|twitter|0.4019|0.0|0.69|0.31|You have my support vote Hillary https://t.co/UvwDw1mA4b
1carpediem2016|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
RandoDaily|GoodOpinionMan|0.0|0.0|1.0|0.0|"@GoodOpinionMan im starting to think that hillary clinton may never be president, but these folks could be onto something"
JacobEngels|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
JacobEngels|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
rugratfarm|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
MyKindOfCrazyMT|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
MyKindOfCrazyMT|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
MelissaTT2000|LisaToddSutton|0.7626|0.135|0.575|0.29|"@LisaToddSutton @KellyannePolls So even our great Hillary or Sanders can not convince U? Hopefully, eventually U will grow up.  Best to U."
ConservativeVO|conservativevoice|0.0|0.0|1.0|0.0|Shes used to it: Hillary Clinton finishes 2nd behind Donald Trump for Times Person of the Year: By  https://t.co/2BiVBvbdQj #conservative
bassyclass|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
PatriotGeorgia|ZKondos|0.0|0.0|1.0|0.0|"RT @ZKondos: @PatriotGeorgia @PatVPeters McCain, a Hillary/Obama/Soros surrogate must be removed from Chairman of the Armed Services comm"
kerrycashion|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
mausiepup|buzz|-0.7269|0.307|0.693|0.0|RT @buzz: When even the foreign power manipulating you is shocked at your party's lack of principle. https://t.co/4erdcrGxSk https://t.co/8
mausiepup|newsweek|-0.7269|0.307|0.693|0.0|RT @buzz: When even the foreign power manipulating you is shocked at your party's lack of principle. https://t.co/4erdcrGxSk https://t.co/8
donaldbroom|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
scott_stalker2|TerriGreenUSA|-0.3612|0.111|0.889|0.0|"RT @TerriGreenUSA: Hillary was careless with her many cell phones and emails. And this happened under Obama's watch, not under a Republican"
b1e56df9ce6549f|GodandtheBear|0.2584|0.0|0.912|0.088|RT @GodandtheBear: I'm not crazy about Hillary is an understatement as to what I feel towards that psychopath. Him being one doesn't change
TrumpInfidel87|funder|-0.9554|0.541|0.459|0.0|@funder #ButcherOfBenghazi Hillary hired terrorists to kill 4 Americans in 2012. Sold firearms to terrorists. THAT IS TREASON. #HangHillary
Axelrod_EJ|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
Bottone6|jfgroves|0.25|0.073|0.813|0.114|"RT @jfgroves: Wait, the woman who offered blowjobs to vote for Hillary is complaining about sexism in the music industry? Lol. https://t."
Bottone6||0.25|0.073|0.813|0.114|"RT @jfgroves: Wait, the woman who offered blowjobs to vote for Hillary is complaining about sexism in the music industry? Lol. https://t."
charawantschoco|ChiIdhoodRuiner|-0.2323|0.317|0.414|0.269|RT @ChiIdhoodRuiner: this leaked email will destroy Hillary's chances of winning https://t.co/MSIra9rnV9
charawantschoco|twitter|-0.2323|0.317|0.414|0.269|RT @ChiIdhoodRuiner: this leaked email will destroy Hillary's chances of winning https://t.co/MSIra9rnV9
Deb1323|kpoulsen|-0.7367|0.275|0.725|0.0|"RT @kpoulsen: Icymi, the ""not sure"" part is that Russia's goal may have been to defeat Hillary, not support her opponent https://t.co/2ubio"
Deb1323|t|-0.7367|0.275|0.725|0.0|"RT @kpoulsen: Icymi, the ""not sure"" part is that Russia's goal may have been to defeat Hillary, not support her opponent https://t.co/2ubio"
txconservgirl|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
CatsTeaRealLife|WalshFreedom|0.5859|0.0|0.84|0.16|"RT @WalshFreedom: If there was evidence that the Russians helped Hillary win, my fellow conservatives would be yelling for an investigation"
Cronyism4Presid|ifunny|0.0|0.0|1.0|0.0|#hillary #hillaryclinton #election https://t.co/yYaqjdG7pL#iFunny https://t.co/8vmVZHmaLk
mamadoc27|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
mrmarkplum|ReaganCoalition|0.0|0.0|1.0|0.0|RT @ReaganCoalition: REVEALED  The Hillary Aide Who KNEW It Was All Over https://t.co/pBxUGkdoYl
mrmarkplum|fiscalconservatives|0.0|0.0|1.0|0.0|RT @ReaganCoalition: REVEALED  The Hillary Aide Who KNEW It Was All Over https://t.co/pBxUGkdoYl
totallmages|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
museisluse|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
rositaagusti|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
rositaagusti|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
nodems16|ramcatalleyetsy|-0.6369|0.394|0.606|0.0|@ramcatalleyetsy @dcexaminer could be Obama hates Hillary n knows she's nuts
rgreen00|MeetThePress|0.0|0.0|1.0|0.0|RT @MeetThePress: Why would Putin hack the U.S. election? Former U.S. Ambassador to Russia Michael @McFaul has a few ideas. WATCH: https://
rgreen00||0.0|0.0|1.0|0.0|RT @MeetThePress: Why would Putin hack the U.S. election? Former U.S. Ambassador to Russia Michael @McFaul has a few ideas. WATCH: https://
Brotherjohnf|brotherjohnf|-0.7845|0.418|0.582|0.0|"New post: Former US Ambassador Attacks First Amendment, Blames Russia Over Hillarys Loss https://t.co/UQVkgZjUpo"
DonnaVishio|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
SSbridges51|Anncostanza1|0.7825|0.094|0.572|0.334|RT @Anncostanza1: Bye Barrack Obama Hillary Clinton Lost Merry Merry Christmas YAY!!!!! #ChristmasIn3Words Bye Harry Reid https://t.co/6G
SSbridges51|t|0.7825|0.094|0.572|0.334|RT @Anncostanza1: Bye Barrack Obama Hillary Clinton Lost Merry Merry Christmas YAY!!!!! #ChristmasIn3Words Bye Harry Reid https://t.co/6G
betz_carl|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
WamplerJim|Evan_McMullin|0.0|0.0|1.0|0.0|@Evan_McMullin @realDonaldTrump if Russia wanted anyone it was hillary... they own the Clintons. America dodged a bullet
Virgil4Trump|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
Virgil4Trump|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
real8BitGeek|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
real8BitGeek|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
GladstoneLaura|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
GladstoneLaura|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
lindarose524|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
RIchgard|jtLOL|0.0609|0.082|0.828|0.09|RT @jtLOL: I'll put it like this: Comey wouldn't have needed to send that letter if Hillary Clinton hasn't been so lawless and paranoid. ht
loisroy72|realjack_bailey|0.0|0.0|1.0|0.0|"RT @realjack_bailey: #Liberals wanted concrete proof from #FBI on #Hillary emails, but will leap to conclusions on #RussiaFBI and CIA #Su"
marktlacroix|immigrant4trump|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
marktlacroix|twitter|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
sunshinette|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
akrinnatus|YouTube|0.4753|0.0|0.819|0.181|I liked a @YouTube video from @markdice https://t.co/4AyM9RpjF0 Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!
akrinnatus|youtube|0.4753|0.0|0.819|0.181|I liked a @YouTube video from @markdice https://t.co/4AyM9RpjF0 Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!
tigertrollz2|CuffyMeh|-0.3071|0.086|0.914|0.0|"RT @CuffyMeh: Russian hacking is bad enough, but just think if Hillary had run all of her classified email thru an unsecure server. Oh man."
Huxley2525|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
teambernie27001|lhfang|-0.6908|0.251|0.749|0.0|RT @lhfang: This guy works for David Brock as a partisan pro-Hillary media critic. And just makes shit up. https://t.co/l3LVbndNDK
teambernie27001|twitter|-0.6908|0.251|0.749|0.0|RT @lhfang: This guy works for David Brock as a partisan pro-Hillary media critic. And just makes shit up. https://t.co/l3LVbndNDK
blaiseking2|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
blaiseking2|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
AlanBigalblack2|bessbell|0.6948|0.217|0.452|0.33|@bessbell @birbigs poor bess flab so starved for attention cheer up sweety hillary loves you but only hillary  LMAO liberal tears
jarianatori|clintonistaa|0.3612|0.0|0.667|0.333|RT @clintonistaa: cheekbones like hillary https://t.co/j0d6T5MJx3
jarianatori|twitter|0.3612|0.0|0.667|0.333|RT @clintonistaa: cheekbones like hillary https://t.co/j0d6T5MJx3
Cory_1077|NozNewz_com|-0.5319|0.186|0.814|0.0|RT @NozNewz_com: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/OSGmSmxWoO
Cory_1077|linkis|-0.5319|0.186|0.814|0.0|RT @NozNewz_com: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/OSGmSmxWoO
FreeSpiritNight|mitchellvii|0.8619|0.0|0.687|0.313|"RT @mitchellvii: Why do these Libs keep saying, ""Hillary won the popular vote!"" That's like saying, ""But we got the most yards!,"" after los"
MyPupVoted|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
IrishSix1|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
lula_reh|wattgirlpower|0.6351|0.0|0.741|0.259|RT @wattgirlpower: Harvard PROF tells @HillaryClinton 2 go to Supreme Court!!  https://t.co/sijKu4qOmt@marciajuell @TyHyCHI @MDBlanchfi
lula_reh|independent|0.6351|0.0|0.741|0.259|RT @wattgirlpower: Harvard PROF tells @HillaryClinton 2 go to Supreme Court!!  https://t.co/sijKu4qOmt@marciajuell @TyHyCHI @MDBlanchfi
Jefd573|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Nieves_18|NiggaTarzan|-0.2348|0.199|0.657|0.143|RT @NiggaTarzan: Me giving my vote to Hillary so Trump doesn't win https://t.co/O7rlfO5ipp
Nieves_18|vine|-0.2348|0.199|0.657|0.143|RT @NiggaTarzan: Me giving my vote to Hillary so Trump doesn't win https://t.co/O7rlfO5ipp
DrHaque|JudicialWatch|0.0|0.0|1.0|0.0|RT @JudicialWatch: In this country our leaders are bound by the rule of law. Hillary Clinton must be held accountable for her actions.http
Mike_Beacham|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
jgsoma|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
jgsoma|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
RebRod|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
RebRod|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
TimidSkye|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
Lisa_Sage|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
billylockner|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
billylockner|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
shad39|HeyTammyBruce|-0.3818|0.167|0.833|0.0|RT @HeyTammyBruce: Hillary Spent Twice As Much As Trump for Her Losing Campaign https://t.co/zuJ1ecioLN
shad39|tammybruce|-0.3818|0.167|0.833|0.0|RT @HeyTammyBruce: Hillary Spent Twice As Much As Trump for Her Losing Campaign https://t.co/zuJ1ecioLN
dutz_neez|AndrewQuackson|-0.2263|0.147|0.853|0.0|RT @AndrewQuackson: The Spetsnaz made Hillary Clinton forget to Campaign in Michigan
TheborderIzsafe|nytimes|-0.7269|0.379|0.621|0.0|Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/Un7wAKMsNX
RickAndKim30yrs|POTUS|-0.4588|0.15|0.85|0.0|Hi @POTUS Remember when Russian Hacks forced Hillary to wipe her server after served a Subpoena to preserve? https://t.co/ArCY5HXbXJ
RickAndKim30yrs|twitter|-0.4588|0.15|0.85|0.0|Hi @POTUS Remember when Russian Hacks forced Hillary to wipe her server after served a Subpoena to preserve? https://t.co/ArCY5HXbXJ
roqchrisy|The_Last_NewsPa|-0.5319|0.177|0.823|0.0|RT @The_Last_NewsPa: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/8uDBCEpH9v https://t.co/WKKUKNWJ
roqchrisy|truthfeed|-0.5319|0.177|0.823|0.0|RT @The_Last_NewsPa: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/8uDBCEpH9v https://t.co/WKKUKNWJ
LelghannMock|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
Balthier28|MadameWoo69|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
Balthier28|change|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
_edwardmondini_|ntvnyr173|0.0|0.0|1.0|0.0|"@ntvnyr173   Everyone thinks Hillary has all this ""experience"":  would we call Benghazi, Libya, Syria &amp; Russia ""experience"" or fiascos?"
PurpleShoesLA|kurteichenwald|-0.2382|0.22|0.67|0.11|"RT @kurteichenwald: No offense, @chucktodd, but when u say no one was sure Russia behind hack pre-election, shows u need to read more. http"
GiveMeLibertyUS|GaetaSusan|-0.8594|0.399|0.498|0.103|"RT @GaetaSusan: Dems, McCain &amp; Graham STOP spreading FAKE NEWS! Every Country hacked Hillary's Private Server! Blame Russia?? What about bl"
CASuperrunner|Keyster101Rich|0.2023|0.098|0.774|0.128|RT @Keyster101Rich: Jill Stein couldn't do it Hillary couldn't do it so now I'll blame the Russian's so much for a peaceful transition from
Doc_Sparky|TrumpSuperPAC|-0.2003|0.144|0.742|0.113|RT @TrumpSuperPAC: #Hillary supporters lying about Hillary's affair with Putin in which she sold 20% of American Uranium to Russia! https:/
Doc_Sparky||-0.2003|0.144|0.742|0.113|RT @TrumpSuperPAC: #Hillary supporters lying about Hillary's affair with Putin in which she sold 20% of American Uranium to Russia! https:/
budb66|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
ktubbs13|Mediaite|0.0|0.0|1.0|0.0|RT @Mediaite: Former U.S. Ambassador to Russia: Vladimir Putin Wanted 'Revenge' on Hillary Clinton https://t.co/e4Kfd6FfcB (VIDEO) https://
ktubbs13|mediaite|0.0|0.0|1.0|0.0|RT @Mediaite: Former U.S. Ambassador to Russia: Vladimir Putin Wanted 'Revenge' on Hillary Clinton https://t.co/e4Kfd6FfcB (VIDEO) https://
CHOCLABLOVER|KailiJoy|-0.6007|0.176|0.824|0.0|"RT @KailiJoy: And now Hillary, who gave us everything of herself and never got a thank you, gets to go on all the goddamned makeup-free hik"
shaycode|JacobRichardsAZ|-0.4215|0.209|0.683|0.108|"RT @JacobRichardsAZ: Hillary would have been a bad president, and on some level I'm glad she lost. But Donald Trump is a continual embarr"
Swift818|AmberleeWhite|-0.3182|0.184|0.703|0.114|@AmberleeWhite @WalshFreedom @SpeakerRyan And Putin and Exxon agreed that Hillary was a threat to their plutarchy.
Tazmanian5|BeachCity55|0.1027|0.077|0.824|0.099|RT @BeachCity55: Jason Chaffetz Forces FBI To Admit They Hid Evidence For Hillary The Entire Time - https://t.co/J6dCFn9KyP
Tazmanian5|proudcons|0.1027|0.077|0.824|0.099|RT @BeachCity55: Jason Chaffetz Forces FBI To Admit They Hid Evidence For Hillary The Entire Time - https://t.co/J6dCFn9KyP
troypotter27|Tymeeks98|0.4019|0.0|0.863|0.137|"RT @Tymeeks98: @mitchellvii @JohnFromCranber Didn't Mexico try to help Hillary, by having Mexican citizens infiltrate US election process?"
julia_alma|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
summerschwab13|AlexErnst|-0.1027|0.11|0.793|0.097|RT @AlexErnst: found out my pet rabbit is a girl and now i'm suddenly mad that hillary clinton isn't the next president of the united states
cocosbentmind|nnwehby_ahmad|0.0|0.0|1.0|0.0|"@nnwehby_ahmad real journalist &amp; people on the ground have said it for years, it's getting harder to lie about now that Hillary's removed."
smell3roses|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Brialalexi|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
Brialalexi|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
norvilgirl|charliekirk11|0.0|0.0|1.0|0.0|"RT @charliekirk11: New evidence shows Russian hackers changed Hillary's speech to include the words ""deplorable and irredeemable"" #FakeNe"
BarbieKayB|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
t_gee_8|NoHoesGeorge|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
t_gee_8|twitter|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
Paxenterris|thehill|-0.2878|0.102|0.898|0.0|@thehill BREAKING: Rothchilds behind massive voter theft for Hillary. A tiny morsel unearthed in WI &amp; MI so recounts were stopped.
robyoungblood11|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
robyoungblood11|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
johncitysq|"elliottkrista,"|-0.2023|0.179|0.684|0.137|"Do you, @elliottkrista, remember Dems said anyone concerned over election integrity was a ""Threat to Democracy""?https://t.co/5YGayG6K1H"
johncitysq|dailywire|-0.2023|0.179|0.684|0.137|"Do you, @elliottkrista, remember Dems said anyone concerned over election integrity was a ""Threat to Democracy""?https://t.co/5YGayG6K1H"
JHarri60|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
JHarri60|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
volpappaw|manny_ottawa|-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
volpappaw||-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
Arexta|ModernDayZorro|-0.3818|0.157|0.843|0.0|RT @ModernDayZorro: Fox News FBI @Wikileaks just took a dump on hillary clinton: https://t.co/SLqPGbcxeh via @YouTube
Arexta|youtube|-0.3818|0.157|0.843|0.0|RT @ModernDayZorro: Fox News FBI @Wikileaks just took a dump on hillary clinton: https://t.co/SLqPGbcxeh via @YouTube
PJConnolly|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TQRlyhHUye via @Change
PJConnolly|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TQRlyhHUye via @Change
hlmartn|gerfingerpoken2|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
hlmartn|americanthinker|-0.7184|0.3|0.7|0.0|"RT @gerfingerpoken2: 3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 htt"
snduffyrn|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
RonCentrelloJr|DailyCaller|-0.296|0.153|0.744|0.103|@DailyCaller I can understand the anger being left out of Hillary's thank you party...pay the money &amp; don't get the ride...
3Panda3|luchadora41|0.0|0.0|1.0|0.0|RT @luchadora41: Were these same voices calling for Hillary Clinton to divest from the Clinton Foundation or CGI while she was Sec. of Stat
cakeman3|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
DKWilson56|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
DKWilson56|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
GADiA_tx|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
VikkiMorgz|bfraser747|-0.6901|0.222|0.778|0.0|"RT @bfraser747:  ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."" ~ @GovMikeHu"
anastasialie83|twitter|0.2158|0.138|0.733|0.13|"I don't want Hillary to bring down the election.I don't want a trump presidency, either.Most importantly, I don https://t.co/PXIEHNovvU"
RebeccaFaussett|FreedomChild3|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
RebeccaFaussett|t|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
PKellyCom|Change|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/ilY2WgK0KZ via @Change
PKellyCom|change|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/ilY2WgK0KZ via @Change
ModernBullWagyu|FishmanLevine|-0.4939|0.158|0.842|0.0|RT @FishmanLevine: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/LQnGEmVzwU vi
ModernBullWagyu|dailycaller|-0.4939|0.158|0.842|0.0|RT @FishmanLevine: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/LQnGEmVzwU vi
YouKeepTheChang|VegasVictory|-0.4939|0.158|0.842|0.0|RT @VegasVictory: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.co/
YouKeepTheChang|t|-0.4939|0.158|0.842|0.0|RT @VegasVictory: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.co/
CarlaMoulton3|Awaken_the_46|0.0|0.0|1.0|0.0|RT @Awaken_the_46: @FaceTheNation @CarlaMoulton3 What's the endgame? Revote? Hillary/Pence? Any GOP is still a puppet &amp; Hillary will have e
Trojan60|GovtsTheProblem|-0.4019|0.325|0.491|0.185|"RT @GovtsTheProblem: Dear Democrats,The Russians didn't make up Hillary Clinton propaganda to stop Hillary. Please stop. I can't stop laug"
paIepeach|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
rockrexx|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
poppylee53152|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
RanchSurfer999|syqau|-0.128|0.13|0.87|0.0|RT @syqau: Alcoholism has contributed to Hillary Clinton's lowered IQ... https://t.co/dxd7hHyqOl
RanchSurfer999|twitter|-0.128|0.13|0.87|0.0|RT @syqau: Alcoholism has contributed to Hillary Clinton's lowered IQ... https://t.co/dxd7hHyqOl
vmlatina|FreedomChild3|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
vmlatina|t|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
BonnieLCollins3|ConservativeFB|-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
BonnieLCollins3||-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
Collette_AZ|sahouraxo|-0.7003|0.28|0.567|0.153|"RT @sahouraxo: Hillary Clinton says #fakenews puts lives at risk.Yeah, like voting for a war that killed millions of innocents based on l"
craig28069746|loug28|-0.2023|0.079|0.921|0.0|@loug28 @babysgramma @Rae_Cass @Cuckerella Hillary armed lybian rebels who turned out to be ISIS. Obama pulled out of Iraq too fast which
Markperugini1|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
roqchrisy|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
SiberiaCat3|MorriseyWV|0.0|0.165|0.671|0.165|".@MorriseyWV @UrlingTreasurer Hillary plans To Help Coal Workers, Trump Has A Scapegoat. #MoralElectors https://t.co/7MVIwSjW02"
SiberiaCat3|npr|0.0|0.165|0.671|0.165|".@MorriseyWV @UrlingTreasurer Hillary plans To Help Coal Workers, Trump Has A Scapegoat. #MoralElectors https://t.co/7MVIwSjW02"
reeltexas|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
reeltexas|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
JanJohnsonFL|RogerJStoneJr|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
JanJohnsonFL|twitter|-0.6486|0.29|0.71|0.0|RT @RogerJStoneJr: Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
TVJMulhern|KrisParonto|-0.3757|0.237|0.643|0.119|@KrisParonto @HillaryClinton @peterdaou So Hillary didn't mock Trump supporters or blame a video? She didn't have a private server?
FisherBurton|BillyVonElds|-0.296|0.099|0.901|0.0|"@BillyVonElds No, we were there with Obama and Hillary bombing Syria &amp; Libya, fucking over Honduras, and monitoring our phones. Fascism."
bill_nusser|smckeon12|0.8314|0.0|0.672|0.328|@smckeon12 not quite but that's ok hey congrats though to you and Hillary on her second place finish
Katherine022610|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Aquasense_USA|nypost|-0.3818|0.224|0.776|0.0|Hillary Clinton's losing campaign cost a record $1.2B https://t.co/sCTpAlGfPu via @nypost
Aquasense_USA|nypost|-0.3818|0.224|0.776|0.0|Hillary Clinton's losing campaign cost a record $1.2B https://t.co/sCTpAlGfPu via @nypost
Stefanyortiz_|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
LabdogEric|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
Maritza03239786|AlisonSpalding2|0.0|0.0|1.0|0.0|RT @AlisonSpalding2: Brazile also got busted fragrantly breaking the laws and ethic of the land by feeding Hillary debate questions. https:
Bipolarization|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
applegherl|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
tpinklittle|HSJECK1|-0.8442|0.349|0.651|0.0|"RT @HSJECK1: Waiting for WaPo to investigate PizzaGate. If it's Fake News, prove it.  Hillary Clinton attacks 'fake news' https://t.co/xy"
tpinklittle|t|-0.8442|0.349|0.651|0.0|"RT @HSJECK1: Waiting for WaPo to investigate PizzaGate. If it's Fake News, prove it.  Hillary Clinton attacks 'fake news' https://t.co/xy"
nana5greatgrand|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
kathyjgabriel|MadameWoo69|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
kathyjgabriel|change|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
SamRomine3|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
EnvyMeGreatly|RepStevenSmith|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
EnvyMeGreatly|dailycaller|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
Sanjay25_|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
JingleBee|SuperSeth64|-0.25|0.08|0.92|0.0|"RT @SuperSeth64: At the moment, Gary Johnson's votes in Florida would push Hillary ahead of Trump. Don't ever talk to me about a protest vo"
CheriCPat|Change|0.0258|0.0|0.945|0.055|"Read this comment, and sign the petition. You exist to prevent a demagogue from assuming this most im... https://t.co/stsMdB09zy via @Change"
CheriCPat|change|0.0258|0.0|0.945|0.055|"Read this comment, and sign the petition. You exist to prevent a demagogue from assuming this most im... https://t.co/stsMdB09zy via @Change"
SM14420071|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
emdharris|unsavoryagents|0.7506|0.0|0.795|0.205|RT @unsavoryagents: THE DEMOCRATS ARE SO CONCERNED ABOUT RUSSIANS HACKING US BUT DON'T SEEM TO CARE THAT HILLARY HAD A STATE DEPARTMENT SER
exhumetw|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
TXCoach10|DineshDSouza|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
TXCoach10|twitter|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
GoykhmanAlla|slone|-0.565|0.207|0.793|0.0|RT @slone: WHO DIDN'T?????????? The list of people who despise Hillary is very long! https://t.co/H3YZOroavx
GoykhmanAlla|twitter|-0.565|0.207|0.793|0.0|RT @slone: WHO DIDN'T?????????? The list of people who despise Hillary is very long! https://t.co/H3YZOroavx
killjoykittens1|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
realnickcarden|mitchellvii|-0.0772|0.16|0.695|0.144|@mitchellvii Yes Bill. Don't you know they forced Donna Brazile to give Hillary debate questions?
LAGRANDIOSA380|CitizensFedUp|0.2023|0.0|0.872|0.128|"RT @CitizensFedUp: Hillary could have legal right to challenge electoral college system and be next US president, says law professor https:"
jaydiener|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
begonefast|thomascolins91|0.5106|0.0|0.751|0.249|"RT @thomascolins91: CA #VOTEHILLARY San Diego Union-Tribune endorsed Hillary Clinton, paper supported Democrat POTUS ~ 1868"
Skeptic4Reason|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
lrnewton1|VivaLaAmes|0.8395|0.091|0.585|0.324|"RT @VivaLaAmes: Me and my daughter love the ""crying for Hillary"" pics. It's like Christmas when you find a new one! This one's a winner! #R"
It_is_NunyaDB|HAGOODMANAUTHOR|-0.798|0.367|0.542|0.091|"RT @HAGOODMANAUTHOR: If Bernie Sanders wasn't cheated, won the nomination, yet lost to Trump, then DEMOCRATS WOULD BLAME BERNIE. Now blame"
JeffreyGSmith|mediaite|-0.7351|0.292|0.708|0.0|"And Trump denies it. ""Former U.S. Ambassador to Russia: Vladimir Putin Wanted Revenge on Hillary Clinton""  https://t.co/4vdVoJukbp"
CindyMae65|TriciasFamily|0.0|0.0|1.0|0.0|"RT @TriciasFamily: https://t.co/RX0q6Ac1fZ Much of Hillary's campaign money came from foreign donors through money laundering,Direct donati"
CindyMae65|westernjournalism|0.0|0.0|1.0|0.0|"RT @TriciasFamily: https://t.co/RX0q6Ac1fZ Much of Hillary's campaign money came from foreign donors through money laundering,Direct donati"
MlchelleMacken|blaubok|0.47|0.096|0.652|0.252|RT @blaubok: When her election was 98% certain - Hillary assured Trump - the election isn't riggedWhen she lost - the election was rigged
linda_wed1|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
expatblackcat|EvelynWhiteGOP|-0.6166|0.237|0.763|0.0|"RT @EvelynWhiteGOP: WATCH  Hillary Calls For CENSORING Conservatives, Her Plan Is SICK https://t.co/5LMuaUi7Sw https://t.co/yrAQudJEOk"
expatblackcat|angrypatriotmovement|-0.6166|0.237|0.763|0.0|"RT @EvelynWhiteGOP: WATCH  Hillary Calls For CENSORING Conservatives, Her Plan Is SICK https://t.co/5LMuaUi7Sw https://t.co/yrAQudJEOk"
Seeitcanbeblank|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
Seeitcanbeblank||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
staggerlee420|Krisp_y|-0.0059|0.192|0.583|0.225|"RT @Krisp_y: Hillary supporters, as highly hypocritical as you are, please repeat after me: ""Russia didn't rig it, she just lost"" https://t"
staggerlee420||-0.0059|0.192|0.583|0.225|"RT @Krisp_y: Hillary supporters, as highly hypocritical as you are, please repeat after me: ""Russia didn't rig it, she just lost"" https://t"
marcylauren|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: Think bout this: Allied intel servives investigating prez-elect 2 learn if he's Putin stooge in place 2 shatter NATO ht
carwizrd|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Me2S3M|jjmikemike|-0.3182|0.187|0.813|0.0|"RT @jjmikemike: Just a reminder from @CNN, from before Hillary lost. https://t.co/xg0c0XllYJ"
Me2S3M|twitter|-0.3182|0.187|0.813|0.0|"RT @jjmikemike: Just a reminder from @CNN, from before Hillary lost. https://t.co/xg0c0XllYJ"
JaniceTXBlessed|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
MsTrishia|SheWhoVotes|0.0|0.0|1.0|0.0|"RT @SheWhoVotes: 1stand this likely isn't Putin's handiworkafter Hillary entered the race with high favorability, the media systematicall"
CaucasianThings|MissMandi00|-0.34|0.231|0.625|0.144|"@MissMandi00 We didnt need ""disinfo"" to hate Hillary. The truth was enough"
Valeriegromes16|btrwkart|0.0|0.0|1.0|0.0|@btrwkart @kiddle https://t.co/XcETfdmQSr
Valeriegromes16|townhall|0.0|0.0|1.0|0.0|@btrwkart @kiddle https://t.co/XcETfdmQSr
1rdgreenberg|charliekirk11|0.8859|0.109|0.523|0.368|@charliekirk11 Russia has is so good that they were able to fix it so Hillary won popular vote &amp; Trump won EC. MSM is so stupid.
SupaReaper|HumanistReport|-0.6705|0.2|0.8|0.0|"RT @HumanistReport: If Hillary Clinton was ever going to denounce fake news, she should have done it after it made her falsely believe Iraq"
organicsgrow|TEN_GOP|0.0|0.0|1.0|0.0|RT @TEN_GOP: 1 Trump didn't take money from Goldman Sachs. 2 Trump owns them.3 Hillary took money from them.4 They own Hillary.Big dif
elijah_azu|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
ZeroAunbis|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
TMB3000|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Cinema_Goulash|Old_Bern_Kenobi|0.4939|0.0|0.814|0.186|@Old_Bern_Kenobi Hillary pretty much pushed Dems so far right they fell off the cliff. #deadparty
PatriotGeorgia|mobile|-0.2263|0.213|0.787|0.0|Hillary pleads to dismiss lawsuit against her https://t.co/anyaFbCiJe
DTROYW63|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
rctu77|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
Trekeee20|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
GiveMeLibertyUS|LindaSuhler|0.4404|0.0|0.847|0.153|RT @LindaSuhler: A good time to mention Hillary Clinton's REAL link to Russia...#RussianHackingShe transferred our uranium to Putin...FOR
RJDownard|DineshDSouza|0.4767|0.122|0.645|0.233|"@DineshDSouza Hillary won popular vote by wide margin, #LoserTrump may yet squeak through Electoral College as losers Harrison &amp; Bush did"
ksenijapavlovic|PavlovicToday|0.0|0.0|1.0|0.0|RT @PavlovicToday: What is the goal of Russian cyber hack? @realDonaldTrump #RussiaHacking #Russia #MAGA #TrumpTransition #Hillary https://
ksenijapavlovic||0.0|0.0|1.0|0.0|RT @PavlovicToday: What is the goal of Russian cyber hack? @realDonaldTrump #RussiaHacking #Russia #MAGA #TrumpTransition #Hillary https://
Konamali1|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Mexicanpov|twitter|0.0656|0.183|0.625|0.192|"LOL, there is So Much wrong doing there, however, in 90mins of pleading his case to DJT in exchange for no pardon o https://t.co/PYxCU8usXR"
sammy27932003|Old_Bern_Kenobi|-0.7579|0.255|0.745|0.0|RT @Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of fac
dms1013|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: Hillary's secret $2.35M Russian Connection was so crooked, even the #CorruptMedia had to covered it. #UraniumOnehttps://t."
jryangolden|CantHardyWait|0.5106|0.107|0.664|0.229|@CantHardyWait @NateSilver538 imagine if Hillary had never got pneumonia and fainted on 9/11 memorial. She wins and Conway looks like a fool
Luvmymariners|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
Luvmymariners||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
oldgeekgal|slone|-0.565|0.207|0.793|0.0|RT @slone: WHO DIDN'T?????????? The list of people who despise Hillary is very long! https://t.co/H3YZOroavx
oldgeekgal|twitter|-0.565|0.207|0.793|0.0|RT @slone: WHO DIDN'T?????????? The list of people who despise Hillary is very long! https://t.co/H3YZOroavx
NeceyDaB0ss|FrankLuntz|-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
NeceyDaB0ss||-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
jkempcpa|LBTheDemocrat|0.1531|0.0|0.918|0.082|@LBTheDemocrat Conmen close deals by pressing flesh &amp; appealing to emotion. Hillary's binders of solid outlined policy were overmatched.
Col_Connaughton|youtube|0.0|0.0|1.0|0.0|Hillary Clinton Faints Part 2 #HACKINGHILLARY https://t.co/WtBgvBsgmM #hillary #clinton #fainting #supported
ClaudiaDAquin|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
koritoprime|OhNoSheTwitnt|-0.68|0.203|0.797|0.0|RT @OhNoSheTwitnt: [Trump on trial for murdering someone on live TV]Defense attorney: But Hillary's emails!Jury: We find the defendant
puffyka81|Col_Connaughton|-0.296|0.145|0.855|0.0|RT @Col_Connaughton: #HILLARY #THIEVERY: Eyewitness #Clinton Foundation Missing from Haitian Aid https://t.co/m1Wo7pt0Yi #corrupt #haiti
puffyka81|youtube|-0.296|0.145|0.855|0.0|RT @Col_Connaughton: #HILLARY #THIEVERY: Eyewitness #Clinton Foundation Missing from Haitian Aid https://t.co/m1Wo7pt0Yi #corrupt #haiti
farmgurl3|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
HiattDon|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
HiattDon|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
GH_obsession|UnBiasedReportr|0.128|0.0|0.927|0.073|RT @UnBiasedReportr: Legal Means That Can Still Make Hillary Clinton The Next U.S. President #Clinton #CIA #Russia #Trump #ElectoralVote ht
teambernie27001|veggie64_leslie|-0.5574|0.204|0.796|0.0|RT @veggie64_leslie: A delusional story about why Hillary lost that captures the lack of responsibility of Clinton and her followers  http
RogerJStoneJr|twitter|-0.6486|0.325|0.675|0.0|Florida #NeverTrump loser Ray Valdes = Crooked Hillary Clinton. He must be stopped. https://t.co/8Bnu81beCn
jaaay_chapman|NoHoesGeorge|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
jaaay_chapman|twitter|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
da_evilgenuis|PrisonPlanet|-0.7351|0.256|0.744|0.0|"RT @PrisonPlanet: Hillary Clinton is concerned about ""fake news"".This is the same woman who claimed the Benghazi attack happened because"
DancesWithPumas|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
lexi_omalley|NoHoesGeorge|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
lexi_omalley|twitter|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
Facetious_man|reckless_mind|0.0|0.0|1.0|0.0|"RT @reckless_mind: @TIME Half the country did not vote. And of the other half, more voted for Hillary Clinton. Where's their story?"
BurnettCynthia|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
BurnettCynthia||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
bepoem|KatieWagnerFox|0.3818|0.134|0.634|0.231|"RT @KatieWagnerFox: Seth Rich narc'd DNC emails because of cheating in Primary to promote Hillary. #SethRich, ultimate Bernie Bro, RIP. #"
ipod49|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
FisherBurton|BillyVonElds|0.3612|0.123|0.737|0.14|@BillyVonElds Sorry. I had no voice when Obama and Hillary were bombing the shit out of Syria &amp; Libya &amp; pushing a Honduras coup. You're off.
wolverines_dad|RNRMississippi|-0.2263|0.215|0.642|0.143|"RT @RNRMississippi: Russians are Amazing: Set up a private server, rigged the primary, used BleachBit to violate a court order, then made"
articcat018|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
mossprinting|LindaSuhler|0.4404|0.0|0.847|0.153|RT @LindaSuhler: A good time to mention Hillary Clinton's REAL link to Russia...#RussianHackingShe transferred our uranium to Putin...FOR
Trillion3|CNN|0.0|0.0|1.0|0.0|@CNN https://t.co/kRF9EM73lH
Trillion3|thegatewaypundit|0.0|0.0|1.0|0.0|@CNN https://t.co/kRF9EM73lH
ArchAngel_Wayne|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
BayShoreIsHome|peopleCRITICamI|0.7427|0.096|0.502|0.402|"REPORT: Hillary Clinton Couldn't Stop Crying, Blamed Comey and Obama for Her Stunning Loss (VIDEO) @peopleCRITICamI  https://t.co/6jpXf5Vvyi"
BayShoreIsHome|thegatewaypundit|0.7427|0.096|0.502|0.402|"REPORT: Hillary Clinton Couldn't Stop Crying, Blamed Comey and Obama for Her Stunning Loss (VIDEO) @peopleCRITICamI  https://t.co/6jpXf5Vvyi"
psmccusker|Love_The_Donald|0.5562|0.085|0.693|0.223|"RT @Love_The_Donald: IN CASE DEMS NEED REMINDER! BOMBSHELL VIDEO: The NSA, not Russia, HACKED the DNC to Help Derail a Hillary Presidency h"
PhoebeMoore11|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
linzucch|BV|0.0|0.0|1.0|0.0|The misjudgments about voters began with Hillary Clinton's announcement video. https://t.co/YFmL9Vt4qn via @BV
linzucch|bloomberg|0.0|0.0|1.0|0.0|The misjudgments about voters began with Hillary Clinton's announcement video. https://t.co/YFmL9Vt4qn via @BV
forgedbytrials|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
BigDuhie1955|9951jackson|0.0|0.0|1.0|0.0|RT @9951jackson: @BigDuhie1955 obama now joined in on the hacking order Cia to look in to the hacking.hillary should be session first thing
histrionicdjh|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Black_Feather55|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
Black_Feather55|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
GJTIII|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
Ferry_Queen|VegasVictory|0.4019|0.0|0.803|0.197|@VegasVictory Hillary donors were expecting quid pro quo. Not interested in philanthropy.
BonnieLCollins3|SheriffClarke|0.4404|0.0|0.884|0.116|RT @SheriffClarke: This is priceless. I would have paid good money to have been on a conference call hook-up when she made this call. https
sunflareweasley|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
AdamAddict|mobile|0.0|0.0|1.0|0.0|  https://t.co/SnFqicCHKy
crw555|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
lulu742|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
lulu742|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
blaiseking2|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
blaiseking2|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
TuxcedoCat|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
marcylauren|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
Hitome29Nygirl|twitter|0.0|0.0|1.0|0.0|#Hillary https://t.co/2xZdAU5glo
jwalkerbryson|ShirlsAdams|0.6249|0.122|0.563|0.315|"@ShirlsAdams @ClaudiaLamb @seriousfun8309 @ericgarland When Hillary and Bernie supporters fight, Trump and his apparatchiks win."
Wareaglebiol|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
Wareaglebiol|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
Hanksingle|katherinejnowak|0.0772|0.104|0.779|0.117|"RT @katherinejnowak: neera has yet to respond with specific errors the dems + hillary's team made; help her out, fam https://t.co/oVuhu75yDS"
Hanksingle|twitter|0.0772|0.104|0.779|0.117|"RT @katherinejnowak: neera has yet to respond with specific errors the dems + hillary's team made; help her out, fam https://t.co/oVuhu75yDS"
Shalom555222|HeyTammyBruce|0.4404|0.0|0.861|0.139|"RT @HeyTammyBruce: Of course. We've been dealing w ""secret"" CIA report revealed to a Hillary supporting blog (WaPost) by anonymous sources."
PatriciaAHenso1|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
rugratfarm|adjordan|0.0|0.0|1.0|0.0|RT @adjordan: Electoral College Make Hillary Clinton President on December 19 - Sign th... https://t.co/Osqx9rWA1a? #ElectoralCollegePetiti
rugratfarm|change|0.0|0.0|1.0|0.0|RT @adjordan: Electoral College Make Hillary Clinton President on December 19 - Sign th... https://t.co/Osqx9rWA1a? #ElectoralCollegePetiti
ProTrump001|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
Rollin_Stone58|veggie64_leslie|-0.5574|0.204|0.796|0.0|RT @veggie64_leslie: A delusional story about why Hillary lost that captures the lack of responsibility of Clinton and her followers  http
McShar1986|ed_hooley|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
McShar1986|truthfeed|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
ipod49|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: I presume you mean Saudi Arabia funding Hillary to the tune of $25 million?No. THAT is not interference at all. https://t.
ipod49||0.0|0.0|1.0|0.0|RT @steph93065: I presume you mean Saudi Arabia funding Hillary to the tune of $25 million?No. THAT is not interference at all. https://t.
70sBaseball|WalshFreedom|0.915|0.0|0.585|0.415|@WalshFreedom could be left's political Hail Mary but you've bought in 100%.  Very noble; I'm sure Hillary supporters would have done same
Sanjay25_|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
TillmanSensei|manny_ottawa|-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
TillmanSensei||-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
inkedcarpenter|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
mariemc11308417|lhfang|0.743|0.0|0.7|0.3|RT @lhfang: Hillary Clinton as Sec of State created a special division within the agency to promote fracking abroad w/Exxon https://t.co/pA
mariemc11308417|t|0.743|0.0|0.7|0.3|RT @lhfang: Hillary Clinton as Sec of State created a special division within the agency to promote fracking abroad w/Exxon https://t.co/pA
gerfingerpoken2|americanthinker|-0.7184|0.333|0.667|0.0|"3 Strikes, Ur Out Hillary. Multiple investigations of felonies American Thinker https://t.co/PMn9JcWweg #PJNET 999 https://t.co/sgSoZqOKCG"
snap_shot_sue|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
deborahjlundy|Tis4Ta|-0.743|0.221|0.708|0.071|"RT @Tis4Ta: I agree with you, &amp; I am mad as hell with why Hillary is not in jail. did she paid everyone off or have deep secrets on them, w"
Trillion3|thehill|0.0|0.0|1.0|0.0|@thehill https://t.co/kRF9EM73lH https://t.co/KGJDwwIMJg
Trillion3|thegatewaypundit|0.0|0.0|1.0|0.0|@thehill https://t.co/kRF9EM73lH https://t.co/KGJDwwIMJg
ModjajiTen|Portosj81J|0.2263|0.0|0.924|0.076|RT @Portosj81J: If the CIA knew that Russia was behind hacking then why did Obama allow Hillary to use a private server with official secre
rollercams|tribelaw|-0.3182|0.161|0.839|0.0|@tribelaw @JoyAnnReid #paytoplay should count to those that relentlessly screamed at Hillary right?
HSJECK1|washingtonpost|-0.8442|0.378|0.622|0.0|"Waiting for WaPo to investigate PizzaGate. If it's Fake News, prove it.  Hillary Clinton attacks 'fake news' https://t.co/xyFSClUfCi"
theocintric|flyer74|-0.8429|0.335|0.665|0.0|RT @flyer74: MR. FAKE NEWS HIMSELF..........ON THE HILLARY CLINTON FOUNDATION DIVISION OF THE CLINTON CRIME FAMILY PAYROLL....... https://t
theocintric||-0.8429|0.335|0.665|0.0|RT @flyer74: MR. FAKE NEWS HIMSELF..........ON THE HILLARY CLINTON FOUNDATION DIVISION OF THE CLINTON CRIME FAMILY PAYROLL....... https://t
shad39|HeyTammyBruce|0.4404|0.0|0.861|0.139|"RT @HeyTammyBruce: Of course. We've been dealing w ""secret"" CIA report revealed to a Hillary supporting blog (WaPost) by anonymous sources."
Sparblack1213|Ian56789|-0.4588|0.13|0.87|0.0|RT @Ian56789: Remember when Russian Hackers forced Hillary to wipe her server after being served with a Congressional Sub Poena to preserve
Charlamaigne|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
allyssar1|twitter|-0.3774|0.269|0.731|0.0|so Hillary lost twice because of.....the Russians...right....lol https://t.co/72SNiZw8d6
pattyjrobinson|jillybobww|0.3612|0.0|0.912|0.088|RT @jillybobww: It is starting to seem like maybe Hillary's email is the one thing the Russians didn't hack &amp; so we should in fact be askin
Canine_Rights|Miami4Trump|0.368|0.129|0.684|0.187|RT @Miami4Trump: Hillary Is FILLED WITH GLEE Because WaPo Is Pushing Her Delusional Conspiracy Theory About Russia Hacking Our Election  #
TMB3000|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
Millenniumistic|MLCzone|0.7351|0.0|0.772|0.228|"RT @MLCzone: As the male power structure hems and haws, Hillary is still winning the popular vote by massive, historic margins. Madame Pres"
LTone|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
LTone||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
mbiancaruddle|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
mbiancaruddle||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
BoCleo2|vivelafra|-0.8977|0.373|0.627|0.0|"RT @vivelafra: This is very sinister.  What this man is describing is an Electoral College coup to unseat #Trump, no doubt exploited by #Hi"
TheMuseCompels|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
loisroy72|AJDelgado13|0.4939|0.101|0.658|0.241|RT @AJDelgado13: Still confused by this theory.Russia meddled to help Trump... and gave Hillary Clinton the popular vote?
mickeypreps|TrumpSuperPAC|-0.4588|0.167|0.833|0.0|"RT @TrumpSuperPAC: The man who hacked #Hillary's personal emails and is currently in prison gave a statement to the legacy media, but they"
glimester|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
BillyVonElds|FisherBurton|0.0731|0.095|0.797|0.109|@FisherBurton would Hillary have filled the cabinet with billionaires too? Maybe. But she wouldn't have restricted inauguration protests
terrij68|JennMarx66|-0.5472|0.15|0.85|0.0|@JennMarx66 what is your point?!? 2.8 million more voted for Hillary are you disputing that? Because you know it is a FACT
Patrici01435181|gerfingerpoken|0.431|0.0|0.831|0.169|RT @gerfingerpoken: (IBD) Hillary Rodham Nixon - Even He Didn't Destroy The Tapes  - https://t.co/OnpEFahSgW - @IBDeditorials - https://t.c
Patrici01435181|investors|0.431|0.0|0.831|0.169|RT @gerfingerpoken: (IBD) Hillary Rodham Nixon - Even He Didn't Destroy The Tapes  - https://t.co/OnpEFahSgW - @IBDeditorials - https://t.c
DavidTravillia1|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Byrlyne|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
JackAppelbaum|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
JackAppelbaum||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
ILPollster|Thor_Sun|0.0|0.0|1.0|0.0|"@Thor_Sun @EricLiptonNYT @ScottShaneNYT @EricLichtblau 2/2 quotes about WMD long before W was in office, including Biden, Hillary, etc."
wolverines_dad|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
for_kent|Isabellaudet|-0.6486|0.371|0.629|0.0|"@Isabellaudet So because Hillary was ""bad"", trump can do no wrong?"
Fastcars2016|LibertyLivesHer|-0.128|0.107|0.805|0.088|@LibertyLivesHer Hillary sure knows how to burn money. Now wonder the country was left broke when both of them left the White House.
SupaReaper|softwarnet|-0.2732|0.091|0.909|0.0|"RT @softwarnet: ""FBI and CIA""Podesta was warned in 2008 to use encryption, Hillary didn't, DNC didn't, Obama's OPM didn't - those who igno"
akondrake|rtyson82|-0.5423|0.304|0.696|0.0|"RT @rtyson82: Hillary still has bad judgment, I see... https://t.co/SK6YONjN7y"
akondrake|twitter|-0.5423|0.304|0.696|0.0|"RT @rtyson82: Hillary still has bad judgment, I see... https://t.co/SK6YONjN7y"
DerekStice|bessbell|-0.2732|0.124|0.876|0.0|@bessbell  honey u must of forgotten Hillary Clinton's Russian reset keep sipping you Mai Tai and leave the the real work to the big boy's
rgreen00|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
Viatcheslavsos3|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
Viatcheslavsos3|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
aarenwent|ChiIdhoodRuiner|-0.4767|0.255|0.745|0.0|"RT @ChiIdhoodRuiner: Forget Trump and Hillary, this man Gary Johnson has no chill  https://t.co/TiTQFMC2xr"
aarenwent|twitter|-0.4767|0.255|0.745|0.0|"RT @ChiIdhoodRuiner: Forget Trump and Hillary, this man Gary Johnson has no chill  https://t.co/TiTQFMC2xr"
mommydean74|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
stevebartin|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
aolghost|Phonycian|-0.2732|0.197|0.678|0.125|RT @Phonycian: Of course Hamas won that election in Palestine which displeased the US and hillarySo they put sanctions on Gaza to starve
gunsrus7|CDCollector23|-0.3818|0.184|0.816|0.0|@CDCollector23 Hillary selling Russia control of uranium mines bothers me. Obama allowing Iran to have nukes bothers me.
CAROLINEMMOOS|twitter|-0.4767|0.171|0.829|0.0|Every so often I remember that Hillary won't be our next president and I am profoundly sad https://t.co/1aMqieWSMx
pammcbide55|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Hispanics16|redflagnews|-0.4019|0.172|0.828|0.0|"Hillary Clinton Spent $1.2 Billion To Lose Election, Twice What Trump Spent https://t.co/km9U4SGznd https://t.co/zcmtqSvPPs"
surrealintel|YourAnonCentral|-0.1779|0.162|0.664|0.174|@YourAnonCentral @cy_guevara So is this posted by Hillary supporters who want to replace Trump with Corporatist War Monger HRC.
Locksley23|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
grocknroll165|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
boblaf|twitter|0.0|0.0|1.0|0.0|The media are all gathering in the bathroom to hear Hillary's next speech. https://t.co/BaPkpAv9Dl
VickiGP1|twitter|0.4168|0.0|0.783|0.217|Hillary still doesn't have a clue. Arrogance is her middle name. https://t.co/dtt7AJLC8a
ZuzzBuzzman|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
BWSchank|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
bbeaty32|AriaWilsonGOP|-0.5255|0.166|0.834|0.0|RT @AriaWilsonGOP: VIDEO : Rush Limbaughs New Hillary Fake News Hit Piece is BLOWING UP the Internet! https://t.co/3hOtjV1lZT https://t
bbeaty32|truthfeed|-0.5255|0.166|0.834|0.0|RT @AriaWilsonGOP: VIDEO : Rush Limbaughs New Hillary Fake News Hit Piece is BLOWING UP the Internet! https://t.co/3hOtjV1lZT https://t
INVUQT|Miami4Trump|0.368|0.129|0.684|0.187|RT @Miami4Trump: Hillary Is FILLED WITH GLEE Because WaPo Is Pushing Her Delusional Conspiracy Theory About Russia Hacking Our Election  #
rachelhamilton_|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
EmpathyNow|JuddLegum|-0.5106|0.221|0.684|0.095|RT @JuddLegum: 9. The GOPs appetite for a hypothetical scandal involving Hillary Clinton is far greater than an actual scandal involving Vl
piercey_judy|nytimes|-0.7269|0.379|0.621|0.0|Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/Ucm53SB9xA
DrHorseshark|QuinnBx|-0.3182|0.247|0.753|0.0|@QuinnBx @LouDobbs #MyBigPollNot mineAbout real reason Ass-Hillary lost
Crossbearer1956|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
Crossbearer1956|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
KamalShaqi|jack3077822|-0.0516|0.139|0.732|0.13|"RT @jack3077822: @oreillyfactor  CHRIS CHRISTIE SIGNED A LAW AGAINST ""BDS"" MOVEMENT WHO BOYCOTT  ISRAEL.  WHEN GEORGE SOROS BIG SUPPORTER"
carwizrd|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
KathyLangeNovak|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
FisherBurton|AlecMacGillis|-0.0772|0.139|0.736|0.126|@AlecMacGillis @TheDeliMan1 So her private server was irrelevant. It's arrogant of you and other Hillary supporters to think otherwise.
danbrady11209|socalmike_SD|0.0|0.0|1.0|0.0|RT @socalmike_SD: Wikileaks: Hillary Clinton Bragged About Being Invited to Putin's 'Inner Sanctum' https://t.co/UyYrkL9WlO via @BreitbartN
danbrady11209|breitbart|0.0|0.0|1.0|0.0|RT @socalmike_SD: Wikileaks: Hillary Clinton Bragged About Being Invited to Putin's 'Inner Sanctum' https://t.co/UyYrkL9WlO via @BreitbartN
MorgLaMignonne|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Billy7004|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
timodonnell14|Duane106|-0.7003|0.266|0.734|0.0|"RT @Duane106: After She Criticized Hillary, 'Morning Joe' Anchor Says NBC Got a Disturbing Call from Clinton Campaign... https://t.co/q6TiV"
timodonnell14|t|-0.7003|0.266|0.734|0.0|"RT @Duane106: After She Criticized Hillary, 'Morning Joe' Anchor Says NBC Got a Disturbing Call from Clinton Campaign... https://t.co/q6TiV"
TrumpetingTrump|WeNeedTrump|-0.296|0.091|0.909|0.0|"RT @WeNeedTrump: Liberals crack me up when they call Trump ""Putin's puppet"" with no evidence. Yet millions of dollars donated to Hillary is"
pammcbide55|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
RonPyke|sullivanamy|0.0|0.0|1.0|0.0|"RT @sullivanamy: That was Joel Benenson's take at U. Chicago a few wks ago. Headlines all scanned as ""emails,"" or ""just more Hillary corrup"
df_mccutcheon|charliekirk11|-0.5106|0.13|0.87|0.0|RT @charliekirk11: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
ggbootsrock|ali|-0.4404|0.112|0.888|0.0|RT @ali: The media won't point to a single thing Hillary Clinton believes or has done outside of the email scandal that Americans may have
Tokaise|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
BernieOrBustLA|Old_Bern_Kenobi|-0.7579|0.255|0.745|0.0|RT @Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of fac
rouleau1|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
PBG2017|realDonaldTrump|-0.4002|0.236|0.583|0.181|"RT @realDonaldTrump: I thought that @CNN would get better after they failed so badly in their support of Hillary Clinton however, since ele"
tzoannop|SenWarren's|0.4256|0.109|0.615|0.277|"Everyone told her so. EVERYONE. No, she chose to support Hillary, whose vested interests stood against @SenWarren's causes."
JamesRitch1|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
JamesRitch1|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
TheMrsDarcy|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Ohboyboy22|cristinalaila1|0.0|0.0|1.0|0.0|RT @cristinalaila1: MSM is more concerned about unsubstantiated claims of Russia hacking the election than Hillary's maid printing up class
kldreams61|PolitixGal|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
kldreams61|twitter|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
hchdwalker|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
JeremyHimli|shoahnuffin1|0.1576|0.286|0.478|0.235|@shoahnuffin1 I didn't help Hillary. I supported the only candidate fit to be President. You supported your Hillary loving man crush.
lapiors|MonicaConCuba|0.0|0.0|1.0|0.0|RT @MonicaConCuba: Algunas vez dijeron que CNN filtr preguntas debate primarias a Hillary Clinton en 2 ocasiones? #MHCC
mark_rector|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
meganbbrennan|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
PatriotRider|JudicialWatch|0.0|0.0|1.0|0.0|RT @JudicialWatch: In this country our leaders are bound by the rule of law. Hillary Clinton must be held accountable for her actions.http
mikecrooks|charliekirk11|0.0|0.0|1.0|0.0|"RT @charliekirk11: Russia potentially being involved is a big deal, but where was the media when Hillary funded her entire staff with forei"
BonnieLCollins3|CronkiteSays|-0.3818|0.205|0.697|0.098|RT @CronkiteSays: REAL NEWSWe've completed an extensive analysis into why Hillary lost and have determined Hillary caused Hillary to lose
PolarWhut|BushwackCA|-0.8109|0.295|0.705|0.0|"RT @BushwackCA: So if #Russia ""Hacked the US election"" then maybe #Hillary didn't win the popular vote. I would bet Russia would rather dea"
HiPaix|prgarc|-0.8655|0.338|0.662|0.0|RT @prgarc: @samsteinhp you mean the part where Obama admin made Hillary LOSE to be able to fight now? That part? Dumb.
dachsiemoron|twitter|0.0|0.0|1.0|0.0|What did he say about Hillary's? https://t.co/8uHktYC1fx
kschoon4|DavidAFrench|-0.3818|0.12|0.88|0.0|"RT @DavidAFrench: Imagine, Republicans, what you would think after losing a close election, then finding out Russia was interfering on Hill"
robinyngbld|change|-0.296|0.239|0.761|0.0|You Can Stop Trump on December 19 https://t.co/3sxsL4n8fS
neiLmunshi|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
neiLmunshi||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
HeysannaHosanna|RepStevenSmith|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
HeysannaHosanna|dailycaller|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
HelenKaufman11|VermillionRich|-0.2732|0.123|0.877|0.0|RT @VermillionRich: .@TrumpUntamed @WalshFreedom @TheLastRefuge2#Hillary has Russian $$ ties &amp; #FakeNews ignores fact INSIDER info = HRC/
reesworld1|ActionTime|0.0516|0.162|0.669|0.169|RT @ActionTime: Trump Backs Off Campaign Promises Again &amp; Again:Trump Admits His Threat to Lock Up Hillary Was Total Lie #Resist #RT https:
takeitstrait|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
realsmile|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
andrelferreiral|RamonCardoso_7|-0.5267|0.239|0.761|0.0|@RamonCardoso_7 @xicosa no queira comparar. No tem como. S bobo caia na conversa que Hillary seria eleita.
Hillary_Rdz|valtrevy|0.0|0.0|1.0|0.0|@valtrevy ah 15 minutos deee
IRBroadshow|DLin71|0.8911|0.0|0.485|0.515|@DLin71 @rznagle She may not have invented sadness but #Hillary surely perfected it.
kaleyiscooool|c0ttin|0.8402|0.0|0.724|0.276|RT @c0ttin: the best christmas present i could ask for is for the electoral college to vote against election results and elect hillary wow
roqchrisy|pRESIDENT_ALIEN|0.0|0.0|1.0|0.0|RT @pRESIDENT_ALIEN: RUSSIA HACKS US NUKESJulius + Ethel Rosenberg get the electric chair. Bill + Hillary Clinton get $100 million.#Fake
ScottRipem99|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
KarmaKittySays|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
KarmaKittySays|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
deborahjlundy|Tis4Ta|-0.1779|0.182|0.657|0.161|"RT @Tis4Ta: Still no lead in Seth Rich death, he work for the government. They should be looking with a fine tooth comb, But for Hillary ev"
GarnerVicky|GustavoRejivik|0.0|0.0|1.0|0.0|@GustavoRejivik @RozierCarol @MrSrsly @BenJealous @mitchellvii He called Hillary on Goldman Sachs speeches. He appoints them to his cabinet!
IreneRosie|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
SiberiaCat3|marceelias|0.555|0.0|0.753|0.247|Plz Help! @marceelias @robbymook @johnpodesta Fate of World In Your Hands. Act NOW! #AuditTheVote #Recount2016 https://t.co/Rze9f8Zpf0
SiberiaCat3|nymag|0.555|0.0|0.753|0.247|Plz Help! @marceelias @robbymook @johnpodesta Fate of World In Your Hands. Act NOW! #AuditTheVote #Recount2016 https://t.co/Rze9f8Zpf0
_nvbodyy|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
isectss|e001|-0.296|0.115|0.885|0.0|"RT @e001: 2016- Dilma caiu- Bonner caiu- Brad Pitt caiu- Hillary caiuSobrou s o Inter, pq time grande no cai."
wrousfljxvm|JohnEkdahl|0.0|0.0|1.0|0.0|RT @JohnEkdahl: Hillary leaves her server open to hacking. Obama rolls over on his belly for Putin for 8 years.  Somehow this is Republican
bbeaty32|wilber7741|-0.6249|0.251|0.685|0.064|RT @wilber7741: Is Hillary rightBREAKING: Hillary Clinton Called Young Voters F*cking Dumb Just Kidding No She Didnt https://t.co/W4UucRM
bbeaty32|t|-0.6249|0.251|0.685|0.064|RT @wilber7741: Is Hillary rightBREAKING: Hillary Clinton Called Young Voters F*cking Dumb Just Kidding No She Didnt https://t.co/W4UucRM
nana5greatgrand|ActualFlatticus|0.2263|0.206|0.557|0.237|"RT @ActualFlatticus: Yes, also Hillary Clinton avoided the entire state of Wisconsin because there are only racists there.  Looking great f"
Fern0947|KellyannePolls|0.3291|0.163|0.661|0.176|@KellyannePolls @Newsweek No but Angela Merkel may have on behalf of Hillary from her warning to Trump after he won the election.
SupaReaper|Tis4Ta|-0.1779|0.182|0.657|0.161|"RT @Tis4Ta: Still no lead in Seth Rich death, he work for the government. They should be looking with a fine tooth comb, But for Hillary ev"
jhorn041159|charliekirk11|0.0|0.0|1.0|0.0|"RT @charliekirk11: New evidence shows Russian hackers changed Hillary's speech to include the words ""deplorable and irredeemable"" #FakeNe"
techindustry|KaylinWinters2|-0.8271|0.386|0.614|0.0|RT @KaylinWinters2: GOP was willing to prosecute Hillary Clinton for fake scandals &amp; lies but evidence of trump colluding with Russia? Not
thekddiamond|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
penny_veritas|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
saints_53|Dovewoman1|0.2023|0.163|0.579|0.258|@Dovewoman1 @WalshFreedom FBI was just trying to play the poor Hillary card. Sympathy votes.
Ladyshrink222|twitter|0.6249|0.052|0.706|0.242|"Yes, Obama and Hillary want to get back at Putin for outsmarting them over the Uranium deal, like that was hard to https://t.co/v4FnArV5ka"
sassygal56222|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
ty00271972|delta1army|0.0|0.0|1.0|0.0|RT @delta1army: Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!  https://t.co/QtkhVcjuW8 via @YouTube
ty00271972|youtube|0.0|0.0|1.0|0.0|RT @delta1army: Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!  https://t.co/QtkhVcjuW8 via @YouTube
RT_CNN|cnn|0.9042|0.0|0.534|0.466|#news #trump #hillary #election #syria CNN Hero of the Year winner: 'God chose me to help' https://t.co/Z8PepbrfpT https://t.co/KomZ8fpMTa
wkirkm|ThankYouDonald|-0.0056|0.094|0.814|0.093|"RT @ThankYouDonald: If Putin really had endorsed Trump, it would have been a blowout. Hillary would have lost bigger than Mondale &amp; Geraldi"
XMerc45|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
SSNjl|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
hollyoptix|JoeWatchesTV|0.755|0.0|0.682|0.318|@JoeWatchesTV Who do u propose for President? Hillary won pop vote. What's your solution to have a Russian state backed leader?
friskydingos|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
JimbauxsJournal|kylegriffin1|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
JimbauxsJournal|theatlantic|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
raklas|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
bbeaty32|wilber7741|0.5023|0.0|0.683|0.317|RT @wilber7741: Is this true regarding Democrats voters?https://t.co/NOTqZM24Fb
bbeaty32|politistick|0.5023|0.0|0.683|0.317|RT @wilber7741: Is this true regarding Democrats voters?https://t.co/NOTqZM24Fb
RT_CNN|twitter|0.0|0.0|1.0|0.0|#news #trump #hillary #election #syria Venezuelan president called a 'Grinch' after toy seizure https://t.co/1FDfNZNSeq
sicg824|EvaSofii|0.0|0.0|1.0|0.0|"@EvaSofii @leslymill @motorhogman @MajBennett @TeamTrumpAZ who ever made outfits for Michelle Obama,Hillary Clinton should make potato sacks"
shortreddog|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
JuliusGoat|metsfan|-0.25|0.143|0.857|0.0|"@metsfan Republican faithless electors breaking for Hillary is the 389,563,208th most likely scenario."
Kimmerjo64|umpire43|-0.5859|0.137|0.863|0.0|RT @umpire43: Hundreds of thousands of Fraud Hillary votes were foung in Detroit and in Millwaukee and in Philly. Did Russia do that to hel
wolfie_tx|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: @AchaPatricia You didnt read a lot of what I wrote pre-election, did you? Try these:https://t.co/JSN8Liptfchttps://t."
wolfie_tx|t|0.0|0.0|1.0|0.0|"RT @kurteichenwald: @AchaPatricia You didnt read a lot of what I wrote pre-election, did you? Try these:https://t.co/JSN8Liptfchttps://t."
AUFanatic23|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
ElCidius|youtube|0.8402|0.0|0.667|0.333|"WOW! Judge Jeanine Pirro makes way too much sense! Speaks Truth about Hillary Clinton, Barack Obama, Putin!! https://t.co/U95UJYOwDr"
JHiker711|FrankLuntz|-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
JHiker711||-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
1776SaveAmerica|Madonna|-0.8521|0.368|0.632|0.0|".@Madonna complains of being called a whore, yet offered blowjobs for @HillaryClinton votes. Must not be good at it. https://t.co/9wud8vehez"
1776SaveAmerica|nytimes|-0.8521|0.368|0.632|0.0|".@Madonna complains of being called a whore, yet offered blowjobs for @HillaryClinton votes. Must not be good at it. https://t.co/9wud8vehez"
PracticalVoter|cfrey01|-0.0516|0.125|0.759|0.116|Sadly too many Americans poorly informed thus trump promises carried the day &amp; Hillary lacked focus direction @cfrey01 @crazylary51
Millenniumistic|UnBiasedReportr|0.128|0.0|0.927|0.073|RT @UnBiasedReportr: Legal Means That Can Still Make Hillary Clinton The Next U.S. President #Clinton #CIA #Russia #Trump #ElectoralVote ht
LandRover1015|EdSkipper|-0.296|0.158|0.731|0.112|RT @EdSkipper: Thanks for this @WalshFreedom It's a crisis. And you know who had a plan to do something about it: Hillary Clinton.
mejehu67|neontaster|0.0|0.0|1.0|0.0|"RT @neontaster: I just realized that Vanquish predicted the future, except that they thought the president working with the Russians would"
GarthDerby|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
deplorable065|realBissell2|0.1779|0.0|0.892|0.108|@realBissell2 @dimensions3x @TopJimy69 @CdotHOW Hillary and Podesta both were into spirit cooking and pedophilia BS......
WizardOfOzballs|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
galinja|KailiJoy|-0.6007|0.176|0.824|0.0|"RT @KailiJoy: And now Hillary, who gave us everything of herself and never got a thank you, gets to go on all the goddamned makeup-free hik"
stevekloscak|hrtablaze|-0.644|0.226|0.774|0.0|RT @hrtablaze: Remember when wikileaks revealed that Primaries were rigged for Hillary? Are the Russians to blame for that too?https://t
stevekloscak||-0.644|0.226|0.774|0.0|RT @hrtablaze: Remember when wikileaks revealed that Primaries were rigged for Hillary? Are the Russians to blame for that too?https://t
lichmearse|rtyson82|-0.8173|0.298|0.702|0.0|"@rtyson82 @CNN Comey, Jill, Gary, and all white people... How many more scapegoats do they need to cover the piss poor decision w Hillary?"
JamesS020770|realjunsonchan|0.4076|0.133|0.632|0.235|"RT @realjunsonchan: -@KellyannePolls completely rekts Rotten Hillary. Lol. This is how America should be governed, spend less, win more. Ni"
Godndguns|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
shazibnadeem|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Fastcars2016|LibertyLivesHer|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
Fastcars2016|vivaliberty|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
datacrown|twitter|0.368|0.158|0.6|0.242|"And George Cooney hates big money in politics, yet he LOVES Hillary. https://t.co/4ALGI1F5oz"
Busa259|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
JohnnyFiorica|Dbargen|0.1531|0.104|0.766|0.131|"RT @Dbargen: Hillary Lost Thanks to One Word, and It's Not 'Russia' @Tom_Blumer #MAGA #TCOT #LNYHBT #DrainTheSwamp #BuildTheWall https://t."
JohnnyFiorica||0.1531|0.104|0.766|0.131|"RT @Dbargen: Hillary Lost Thanks to One Word, and It's Not 'Russia' @Tom_Blumer #MAGA #TCOT #LNYHBT #DrainTheSwamp #BuildTheWall https://t."
tariq_alauddin|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
TinaDuryea|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
ilrahmawat1|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
ilrahmawat1|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
Anyshka|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
Mc_Heckin_Duff|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
cassidyphoenyx|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
cassidyphoenyx|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
Nohillary2|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
flyer74|flyer74|0.0|0.0|1.0|0.0|RT @flyer74: THIS BOOK IS BEING WRITTEN BY HILLARY CLINTON https://t.co/tQJyoJvgQY
flyer74|twitter|0.0|0.0|1.0|0.0|RT @flyer74: THIS BOOK IS BEING WRITTEN BY HILLARY CLINTON https://t.co/tQJyoJvgQY
beatlebabe49|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
KarmaKittySays|nia4_trump|-0.7184|0.304|0.696|0.0|"RT @nia4_trump: #FridayFeeling Hillary emerged 3 times since her crushing defeat, always wearing purple, the color of Rebellion &amp; Power.  V"
jamien8926|qstafford50|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
jamien8926|palmerreport|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
RCakora|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
RCakora|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
JohnBlast2000|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
Kyriati|good|0.3774|0.0|0.861|0.139|"The icon for the Rock if you pick female is Hillary Clinton, so thats cool https://t.co/8j21e8IIxN https://t.co/kCIHAuSsdP"
ConsiderThis1|silvanet|-0.5859|0.275|0.725|0.0|Hillary's Primary Election Fraud is the FORCING I was talking about. @silvanet
RealJimPeterson|CarmineZozzora|0.85|0.0|0.634|0.366|RT @CarmineZozzora: Russian hacking narrative mysteriously absent when Hillary was sure to win - but magically surfaces after Trump's win?
Maggieknp|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
mj_schwarz|BobMcElvaine|0.5574|0.0|0.816|0.184|RT @BobMcElvaine: Hillary Can Be a Hero by Saving America from Trump https://t.co/J6H79uNWGv via @HuffPostPol #Hillary #StopTrump #Electora
mj_schwarz|huffingtonpost|0.5574|0.0|0.816|0.184|RT @BobMcElvaine: Hillary Can Be a Hero by Saving America from Trump https://t.co/J6H79uNWGv via @HuffPostPol #Hillary #StopTrump #Electora
KarmaKittySays|BrittPettibone|0.4404|0.0|0.861|0.139|"RT @BrittPettibone: #ImStillNotOver the fact that, based on zero evidence, Hillary Supporters insist that Russian Hackers interfered in the"
deanawa55339161|TriciasFamily|0.0|0.0|1.0|0.0|"RT @TriciasFamily: https://t.co/RX0q6Ac1fZ Much of Hillary's campaign money came from foreign donors through money laundering,Direct donati"
deanawa55339161|westernjournalism|0.0|0.0|1.0|0.0|"RT @TriciasFamily: https://t.co/RX0q6Ac1fZ Much of Hillary's campaign money came from foreign donors through money laundering,Direct donati"
exhumetw|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
NightShiftNews|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
NightShiftNews|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
xpro1|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
NYlovesTrump|An0nKn0wledge|-0.6739|0.171|0.829|0.0|RT @An0nKn0wledge: THERE IS MORE EVIDENCE OF ALIENS EXISTING THEN THE RUSSIANS HACKING THE ELECTION.. BTW THE ELECTION FRAUD SO FAR ALL IN
bzazzie|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: #PodestaEmails more proof of Hillary's Russian Connections. ""Grassley Letter"" to Loretta Lynch. #CorruptMedia let this stor"
goldcamaro|ladygaga|-0.4404|0.139|0.861|0.0|RT @ladygaga: If you feel scared about the current state of American politics and Whitehouse sign this petition: https://t.co/2K88hLD8hn
goldcamaro|change|-0.4404|0.139|0.861|0.0|RT @ladygaga: If you feel scared about the current state of American politics and Whitehouse sign this petition: https://t.co/2K88hLD8hn
gc_cic|TrinityNYC|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
gc_cic|t|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
CocoThePatriot|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
JeffersonsNotes|westernlvr|-0.5994|0.353|0.647|0.0|"@westernlvr Had Russia made Hillary president, no problem? I don't think so."
csluna1ruby|intlspectator|0.8689|0.0|0.634|0.366|"RT @intlspectator: Hillary Clinton's popular vote lead now at 2.8 million votes, the greatest popular vote victory for presidential electio"
USAHipster|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
FaithfulChickie|ClutchScience|0.7777|0.0|0.726|0.274|@ClutchScience Hillary wasn't the runner-up! She won by 2.7 mil. votes.In a true democracy the person w/most votes is the winner.@ezlusztig
mlw975|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
YouKeepTheChang|TheSantaParty|-0.4939|0.167|0.833|0.0|RT @TheSantaParty: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - https://t.co/jALmHrnlkL
YouKeepTheChang|vivaliberty|-0.4939|0.167|0.833|0.0|RT @TheSantaParty: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - https://t.co/jALmHrnlkL
bsdesigns18|conservativetribune|-0.4472|0.283|0.575|0.142|"Hillary Whines About Fake News, So Rush Runs Special 90-Second Montage Just for Her https://t.co/x4m5BrrPXk"
rharrisonfries|slone|-0.4466|0.118|0.882|0.0|RT @slone: We KNOW that McCain and Graham voted for Hillary b/c they're both GLOBALISTS. There is NO difference btwn a D globalist &amp; an R g
chidiebereogbe1|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
chidiebereogbe1|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
_royallytatoox|HillaryTheBOSS|0.0|0.0|1.0|0.0|RT @HillaryTheBOSS: Hillary del Rodman  https://t.co/O5aanBZoQd
_royallytatoox|twitter|0.0|0.0|1.0|0.0|RT @HillaryTheBOSS: Hillary del Rodman  https://t.co/O5aanBZoQd
904Activist|truthrevolt|0.0|0.0|1.0|0.0|https://t.co/Mprcse6wuR https://t.co/RIjVGJy4D4
exhumetw|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
parklochu|maItinerecords|0.4019|0.0|0.838|0.162|RT @maItinerecords: hillary clinton flew all the way to hong kong to support twice https://t.co/Dsmufj6Xes
parklochu|twitter|0.4019|0.0|0.838|0.162|RT @maItinerecords: hillary clinton flew all the way to hong kong to support twice https://t.co/Dsmufj6Xes
chenoehart|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
ElisaMichaels|twitter|-0.7717|0.261|0.739|0.0|".Too late. #Obama knew #Hillary had a private server in violation of law. He's an accomplice to crime, if not compl https://t.co/v4Otj3ogfV"
patty_restaino|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
meow2u22|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
deborahjlundy|Old_Bern_Kenobi|-0.7579|0.255|0.745|0.0|RT @Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of fac
GraysonBlount|WhitePeepsDo|-0.4767|0.255|0.745|0.0|"RT @WhitePeepsDo: Forget Trump and Hillary, this man Gary Johnson has no chill https://t.co/c5nOgggTd8"
GraysonBlount|twitter|-0.4767|0.255|0.745|0.0|"RT @WhitePeepsDo: Forget Trump and Hillary, this man Gary Johnson has no chill https://t.co/c5nOgggTd8"
crebj|TheTakeaway|-0.2023|0.239|0.556|0.205|"@TheTakeaway @PRI @WNYC Hillary Clinton. She's no loser, is a graceful conceder, and would have been a fine president."
SJSciarra|JuddLegum|0.0|0.0|1.0|0.0|RT @JuddLegum: 1. Let's go back to Hillary's email server for a minute. What was the concern?
RoselaMetal|Change|0.0|0.0|1.0|0.0| Sign the Petition!  Electoral College: Make Hillary Clinton President on December 19  https://t.co/L60zpgh8Bu https://t.co/iR0TxMoPmK
capricorniall|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
JtMobleyFla|HillaryClinton|-0.2732|0.155|0.744|0.101|"THE LEAK IS USA,DNI, DHS THAT DID NOT WANT @HillaryClinton their boss, deal with it Hillary https://t.co/MUQgguXaX3"
JtMobleyFla|twitter|-0.2732|0.155|0.744|0.101|"THE LEAK IS USA,DNI, DHS THAT DID NOT WANT @HillaryClinton their boss, deal with it Hillary https://t.co/MUQgguXaX3"
Rosechristenbe1|Peterthegreat16|0.1027|0.13|0.688|0.181|"RT @Peterthegreat16: @TPH_news @realDonaldTrump hillary won 57 out of 3,143 counties. Who gives a shit what LA and NYC want. They don't rep"
rebfansr|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
mowser1970|CarmineZozzora|-0.7906|0.269|0.731|0.0|RT @CarmineZozzora: The FBI that covered for Hillary's serial felonies to conceal her past felonies is protecting Donald Trump now?Got fa
exhumetw|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: The Democrats all debate who's going to get out of Hillary's way first, except for VERMONT'S OWN BERNIE SANDERS, who...get"
rgreen00|bfraser747|-0.6901|0.222|0.778|0.0|"RT @bfraser747:  ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."" ~ @GovMikeHu"
Deemoney521|janet_yackle|-0.3612|0.167|0.739|0.094|"RT @janet_yackle: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/MoUSXY0OP6 via @crooksandlia"
Deemoney521|crooksandliars|-0.3612|0.167|0.739|0.094|"RT @janet_yackle: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/MoUSXY0OP6 via @crooksandlia"
RealtorBo|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
RealtorBo|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
allofusfortrump|bfraser747|-0.6901|0.222|0.778|0.0|"RT @bfraser747:  ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."" ~ @GovMikeHu"
seedcollector|andersonDrLJA|-0.7783|0.31|0.596|0.094|"RT @andersonDrLJA: UNBELIEVABLE LIBERAL LOGIC!!!#HILLARY LOSES BIG TIME WITH BIG FACTOR BEING HER CRIMINAL BEHAVIOR!  THEN, SHE &amp; LIBERAL"
hale4jesus|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
CROWENATION2016|RepStevenSmith|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
CROWENATION2016|dailycaller|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
Tuscan21_PM|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
_corpp|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
_corpp|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
DKWilson56|sullivanamy|0.0|0.0|1.0|0.0|"RT @sullivanamy: That was Joel Benenson's take at U. Chicago a few wks ago. Headlines all scanned as ""emails,"" or ""just more Hillary corrup"
MLCzone|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
LaurieRobert6|greggutfeld|-0.2528|0.246|0.594|0.16|"@greggutfeld @GregGutfeldShow Scandal. Hillary dilarry flock, bickering won't stop."
lionking_007|2ALAW|-0.3182|0.223|0.777|0.0|RT @2ALAW: @LeahR77 @SenJohnMcCain @LindseyGrahamSC Hillary Sees A Ghost https://t.co/EOvIdoE4iU
lionking_007|twitter|-0.3182|0.223|0.777|0.0|RT @2ALAW: @LeahR77 @SenJohnMcCain @LindseyGrahamSC Hillary Sees A Ghost https://t.co/EOvIdoE4iU
tobyonekonobe|BurtEichenwald|-0.1531|0.086|0.914|0.0|"RT @BurtEichenwald: @mtracey @BillMoranWrites And then, without any facts, saying it affected the 4 closest states and Hillary otherwise"
SolarGuacha|TrumpSuperPAC|-0.4588|0.167|0.833|0.0|"RT @TrumpSuperPAC: The man who hacked #Hillary's personal emails and is currently in prison gave a statement to the legacy media, but they"
cdsmith42|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
Clay_Scott_|owasow|0.0|0.348|0.303|0.348|@owasow truth: Hillary lost
Manchu71|CholericCleric|0.462|0.073|0.772|0.155|@CholericCleric I dislike Fox but why give it so much credit? Liberal rags descended to Sanjay Jha level pompom waving for Hillary
toby1995|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
UWantMyVote_Why|atleecs|0.1406|0.082|0.816|0.102|@atleecs @SenatorBoxer Maybe Hillary's being quiet &amp; letting this play out. Then Trump has no reason 2 go after her &amp; take focus off himself
trillcyberdad|twitter|0.0|0.0|1.0|0.0|didn't he also vow to investigate hillary? https://t.co/JHgT6UTXEi
2Twitte39301335|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
2Twitte39301335|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
cfknnyc|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
AlPal_Lehman|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
amerycarlson|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
carolina_brenna|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
RalphHornsby|thegatewaypundit|0.2732|0.132|0.683|0.185|Hillary Clinton Spent $1.2 Billion to Lose Election - TRUMP Spent Around $600 Million to Win https://t.co/oECrCYEYXJ
nancydmoore25|DineshDSouza|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
nancydmoore25|twitter|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
snowstorm1944|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Col_Connaughton|youtube|-0.296|0.167|0.833|0.0|#HILLARY #THIEVERY: Eyewitness #Clinton Foundation Missing from Haitian Aid https://t.co/m1Wo7pt0Yi #corrupt #haiti
AngelicPrado|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
AngelicPrado|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
Nottinghams1|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
Nottinghams1|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
xrfauxtard|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
Landry777Tom|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
hartfordwolf|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
NatashaLifecoac|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
artblam|dailymail|0.0|0.0|1.0|0.0|Hillary is confirmed KGB. Clinton says she'd rather have dinner with Putin than Trump https://t.co/kpkFQfserq https://t.co/oQ0ZNi4Jm4
OddLane|reason|0.0|0.0|1.0|0.0|The First Amendment as suggestion box: https://t.co/jQ45zepGyP #HillaryClinton #Fakenews
jebanamac|DSORennie|0.0|0.0|1.0|0.0|@DSORennie Talk about Foreign influence. Did Russian hackers force Hillary to take millions in Saudi money?
valtrevy|Hillary_Rdz|0.0|0.0|1.0|0.0|@Hillary_Rdz jajaja en San Nico
hnvance40|SharonMcCutchan|-0.4939|0.167|0.833|0.0|RT @SharonMcCutchan: Senator D'Amato Drops Bomb: Hillary Allowed Russia to Take Ownership of ... https://t.co/kVjS4EYc9O via @YouTube
hnvance40|youtube|-0.4939|0.167|0.833|0.0|RT @SharonMcCutchan: Senator D'Amato Drops Bomb: Hillary Allowed Russia to Take Ownership of ... https://t.co/kVjS4EYc9O via @YouTube
Sheilahoover12|umpire43|0.0|0.0|1.0|0.0|RT @umpire43: In Millwaukee day 5 of recount Hillary had 356000 votes thrown out for Fraud.Boxes in Millwaukee did not match poll books RUS
Anyshka|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
stillval13|arunanaimji|0.644|0.0|0.701|0.299|@arunanaimji @FoxNews @foxnewspolitics and who do you trust? Hillary? Bernie? Jill?
Maimaimaire|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
boggs_69|Uberpatroit|-0.296|0.121|0.879|0.0|@Uberpatroit @Billhic02785574 @NateSilver538 And Saddam had WMD's....you Hillary sychophants are priceless...now the CIA can do no wrong...
martucci_peter|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
validthought|AlphaHuskyAlpha|0.4973|0.0|0.801|0.199|@AlphaHuskyAlpha @NickNoelte1 Did Hillary have secret meetings with intl bankers? Yup. Facts aren't racist.
oceandog|nypost|-0.3818|0.224|0.776|0.0|Hillary Clinton's losing campaign cost a record $1.2B https://t.co/EklVFrpHsG via @nypost
oceandog|nypost|-0.3818|0.224|0.776|0.0|Hillary Clinton's losing campaign cost a record $1.2B https://t.co/EklVFrpHsG via @nypost
SiberiaCat3|walterbegayjr|0.4926|0.0|0.814|0.186|.@walterbegayjr @robertsgraham Hillary has a better tax plan. Don't Vote Trump he's for himself! #MoralElectors https://t.co/N8jmYpCLYI
SiberiaCat3|youtube|0.4926|0.0|0.814|0.186|.@walterbegayjr @robertsgraham Hillary has a better tax plan. Don't Vote Trump he's for himself! #MoralElectors https://t.co/N8jmYpCLYI
AnacVentilari|America_1st_|-0.3612|0.143|0.857|0.0|"RT @America_1st_: Reince Priebus: ""The Russians didnt tell Hillary Clinton to ignore Wisconsin or Michigan."" https://t.co/xkRn0HnAh4"
AnacVentilari|twitter|-0.3612|0.143|0.857|0.0|"RT @America_1st_: Reince Priebus: ""The Russians didnt tell Hillary Clinton to ignore Wisconsin or Michigan."" https://t.co/xkRn0HnAh4"
KarmaKittySays|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
ModjajiTen|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
MarkChesney|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
YReag|AIIAmericanGirI|0.5411|0.0|0.741|0.259|@AIIAmericanGirI Russia hired Huma Abedin has the right hand to Hillary!
AlisaaGail|HumanistReport|-0.6705|0.2|0.8|0.0|"RT @HumanistReport: If Hillary Clinton was ever going to denounce fake news, she should have done it after it made her falsely believe Iraq"
tobyonekonobe|veggie64_leslie|0.2584|0.0|0.873|0.127|RT @veggie64_leslie: @mtracey @soso_koba @NateSilver538 Especially when he knew Hillary didn't bother to campaign https://t.co/q1wzXr8674
tobyonekonobe|twitter|0.2584|0.0|0.873|0.127|RT @veggie64_leslie: @mtracey @soso_koba @NateSilver538 Especially when he knew Hillary didn't bother to campaign https://t.co/q1wzXr8674
ArtCareServices|GeorgeShiber|0.0|0.0|1.0|0.0|RT @GeorgeShiber: Tell me again exactly what Hillary did wrong?! With all the 'external forces' and she still beat every man in history: 'g
TheMissWare|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
joselinda69|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
FidTradZ101|SugarspotAnnie|0.6369|0.0|0.811|0.189|"@SugarspotAnnie @Adsocheetie @beulahcrusoe @patticakeski @PenPure1  Hillary was all for that, tried to do it here. But socialists love her."
Fastcars2016|eSeSthetics|-0.5267|0.195|0.805|0.0|@eSeSthetics @paulmeyer745 @Cantkillrspirit @trump2016fan @TAGOS22 To puke on their faces; Esp on Hillary's and G.Soros. 
PavlovicToday|realDonaldTrump|0.0|0.0|1.0|0.0|What is the goal of Russian cyber hack? @realDonaldTrump #RussiaHacking #Russia #MAGA #TrumpTransition #Hillary https://t.co/Cl8nXv99Ql
PavlovicToday|twitter|0.0|0.0|1.0|0.0|What is the goal of Russian cyber hack? @realDonaldTrump #RussiaHacking #Russia #MAGA #TrumpTransition #Hillary https://t.co/Cl8nXv99Ql
Curtlando|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
RyanResign|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
SallyJupiterRA|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
SallyJupiterRA||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
CocoThePatriot|tteegar|-0.3182|0.095|0.905|0.0|RT @tteegar: .@PrisonPlanet Libtards b likeHow many ways can we rub a historic Hillary Clinton loss in &amp; pour salt on this wound we con
IrishSix1|DaysOfTrump|-0.5994|0.196|0.804|0.0|"RT @DaysOfTrump: #AmericaFirst Patriots inside USgov are waging a civil war w international socialists (Hillary, Soros..) that have infiltr"
Natalydubai|RepStevenSmith|0.0772|0.0|0.939|0.061|RT @RepStevenSmith: Want to hear about what Hillary did in Libya from a real journalist? @wikileaks Julian Assange explains it in 2 minutes
mikew6161|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
coniinthegarden|ProgressiveArmy|-0.2263|0.128|0.872|0.0|Donald Hasnt Forgotten About Hillarys Emails and Neither Have House Republicans https://t.co/9BTGMPMZaV via @ProgressiveArmy
coniinthegarden|progressivearmy|-0.2263|0.128|0.872|0.0|Donald Hasnt Forgotten About Hillarys Emails and Neither Have House Republicans https://t.co/9BTGMPMZaV via @ProgressiveArmy
StormSpinning|AdamParkhomenko|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
StormSpinning|nydailynews|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
Proud4USA1|dongsmack|0.3612|0.0|0.839|0.161|Thank U Rock ( @dongsmack ) for coming forward 2 prove Hillary is right. Deplorable misogynists exist. https://t.co/zmBO2ZfE0y
Proud4USA1|twitter|0.3612|0.0|0.839|0.161|Thank U Rock ( @dongsmack ) for coming forward 2 prove Hillary is right. Deplorable misogynists exist. https://t.co/zmBO2ZfE0y
yanson07230606|TrinityNYC|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
yanson07230606|t|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
LogjamminPete|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
purpledalmation|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
purpledalmation|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
braunaa|danpfeiffer|-0.7096|0.277|0.723|0.0|RT @danpfeiffer: I am confused. Were voters supposed to takes Trump's attacks on Hillary's ties to Goldman Sachs literally or seriously? ht
kolnhausen|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
cosmogenesis777|worldnewsdailyreport|0.0|0.0|1.0|0.0|"Yoko Ono: ""I Had an Affair with Hillary Clinton in the '70s"" https://t.co/Zxd3c3HNmt"
dmneedham|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
MyPlace4U|LVNancy|0.5719|0.0|0.791|0.209|"RT @LVNancy: #RussianHackers IF sore-Loser, Hillary had won, would we be having this conversation?#SundayMorning #TRUMP#AmericaFirst"
dlreinbeau|Krisp_y|-0.0059|0.192|0.583|0.225|"RT @Krisp_y: Hillary supporters, as highly hypocritical as you are, please repeat after me: ""Russia didn't rig it, she just lost"" https://t"
dlreinbeau||-0.0059|0.192|0.583|0.225|"RT @Krisp_y: Hillary supporters, as highly hypocritical as you are, please repeat after me: ""Russia didn't rig it, she just lost"" https://t"
stp_han|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
AmericanMom2|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
sherrysue66|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
sarahsettgo|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
womenaresmarter|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
Hrgrthr71|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
h0memadetweets|twitter|-0.6124|0.406|0.438|0.156|Defeating Hillary Clinton feels like a war victory. #AmericaisBack #MAGA https://t.co/AZYPPGFXmu
Stormysu|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
counting76cou|S1776frdm|-0.9186|0.519|0.417|0.064|"RT @S1776frdm: Hillary Sucked at everything except Treason Corruption Pay4PlayKindness of Spirit Racism, Hate 4 Average Citizens--https:/"
counting76cou||-0.9186|0.519|0.417|0.064|"RT @S1776frdm: Hillary Sucked at everything except Treason Corruption Pay4PlayKindness of Spirit Racism, Hate 4 Average Citizens--https:/"
GiuseppeSab|DailyCaller|-0.8126|0.359|0.641|0.0|RT @DailyCaller: Shooting The Wrong Messenger  Morning Joe Calls Out Hillary Clinton For Hiding Behind Fake News https://t.co/gq71mB
GiuseppeSab|t|-0.8126|0.359|0.641|0.0|RT @DailyCaller: Shooting The Wrong Messenger  Morning Joe Calls Out Hillary Clinton For Hiding Behind Fake News https://t.co/gq71mB
mosfoodographer|nypost|-0.5106|0.452|0.548|0.0|@nypost @realDonaldTrump Hillary for Prison
anastasiakhramo|twitter|-0.2755|0.19|0.81|0.0|Because they don't like Hillary Clinton? Durgh. Face palm. https://t.co/pYYkCXE7RS
BubbaLiberal|briantashman|0.4767|0.0|0.846|0.154|RT @briantashman: Donald Trump doesn't listen to the intelligence community. But he does listen to this guy https://t.co/Er5TdMuPEn
BubbaLiberal|rightwingwatch|0.4767|0.0|0.846|0.154|RT @briantashman: Donald Trump doesn't listen to the intelligence community. But he does listen to this guy https://t.co/Er5TdMuPEn
slowbob|YouTube|0.0|0.0|1.0|0.0|Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!  https://t.co/CW9wj3kqBa via @YouTube
slowbob|youtube|0.0|0.0|1.0|0.0|Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!  https://t.co/CW9wj3kqBa via @YouTube
Brendag38323989|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
joecuts134|TroyCoby|0.0|0.0|1.0|0.0|RT @TroyCoby: Hillary Clinton has been drinking a lot... https://t.co/vPJh1ZkOFN
joecuts134|twitter|0.0|0.0|1.0|0.0|RT @TroyCoby: Hillary Clinton has been drinking a lot... https://t.co/vPJh1ZkOFN
ValiantSentry|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
ValiantSentry|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
DAndalora_Bella|ThinkCenter1968|-0.5267|0.129|0.871|0.0|RT @ThinkCenter1968: This was actually announced at some point back in the campaign so it seems Hillary &amp; Obama R openly lying about the ma
princesskimcj|ArianeBellamar|0.5719|0.0|0.837|0.163|"RT @ArianeBellamar: @realDonaldTrump  Hillary won EVERY major economy in EVERY state, proving that the most under-educated ppl in this co"
gilberthoughton|WhitePeopIeCray|0.0|0.0|1.0|0.0|"RT @WhitePeopIeCray: ""Hillary for prison!!""""Let's make it happen"" https://t.co/TuNeWBefoB"
gilberthoughton|vine|0.0|0.0|1.0|0.0|"RT @WhitePeopIeCray: ""Hillary for prison!!""""Let's make it happen"" https://t.co/TuNeWBefoB"
DAILYBLUEblog|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
roqchrisy|Democrat_4Trump|0.3182|0.116|0.667|0.218|RT @Democrat_4Trump: Hillary Clinton's losing campaign cost a record $1.2B and MANY LIVES of innocent people like Seth. https://t.co/hLCoph
roqchrisy|t|0.3182|0.116|0.667|0.218|RT @Democrat_4Trump: Hillary Clinton's losing campaign cost a record $1.2B and MANY LIVES of innocent people like Seth. https://t.co/hLCoph
Just_A_Bill_|liars_never_win|-0.5423|0.171|0.829|0.0|RT @liars_never_win: It wasn't the hacking of Podesta's emails that made Hillary look bad. It was the content
luvmom8702|JSavoly|0.2263|0.0|0.872|0.128|"RT @JSavoly: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton #StollenElection #ComradeTrump  https://t.co/LyFMVe3WP0"
luvmom8702|crooksandliars|0.2263|0.0|0.872|0.128|"RT @JSavoly: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton #StollenElection #ComradeTrump  https://t.co/LyFMVe3WP0"
geokaren|twitter|0.5423|0.0|0.759|0.241|Putin just wants power and control. Hillary was an added bonus. https://t.co/8s3SNbUhPs
De5p|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
De5p|t|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
KOMBUCHABABY|Old_Bern_Kenobi|-0.7579|0.255|0.745|0.0|RT @Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of fac
HelenKaufman11|PolitixGal|0.0|0.0|1.0|0.0|RT @PolitixGal: THE REAL HILLARY... https://t.co/MYCYvoXy3B
HelenKaufman11|twitter|0.0|0.0|1.0|0.0|RT @PolitixGal: THE REAL HILLARY... https://t.co/MYCYvoXy3B
Tortured_Verse|PaulDeCampo|0.4019|0.0|0.856|0.144|"@PaulDeCampo I was taunting @one110731 about alleged ""leftists"" in USA. Hillary &amp; Democrats are center-left. Definitely not ""leftists."""
CheeperSteeper|Hispanics16|-0.4767|0.171|0.829|0.0|"RT @Hispanics16: Joe Scarborough: HILLARY CLINTON COST HILLARY CLINTON THE ELECTION, Not Fake News https://t.co/vaw8FwlP1r https://t.co/j"
CheeperSteeper|usapoliticstoday|-0.4767|0.171|0.829|0.0|"RT @Hispanics16: Joe Scarborough: HILLARY CLINTON COST HILLARY CLINTON THE ELECTION, Not Fake News https://t.co/vaw8FwlP1r https://t.co/j"
kc6ymp|TheRealN6BHU|-0.5267|0.152|0.848|0.0|@TheRealN6BHU @MotherJones it's a conspiracy uncle Donnie is going after all the pantie waving Hillary liberals OMG that's you right Dave 
hyland114|twitter|-0.875|0.417|0.583|0.0|"FAKE NEWS GUY CHUCK TODD, NEVER QUESTIONED HILLARY ABT CLASSIFIED EMAIL FIASCO N CLASSIFIED INFO HACK. BENGHAZI, https://t.co/QLEMIx2Qon"
DanielAPfister|patrickhealynyt|0.8519|0.0|0.491|0.509|Great feature on Madonna &amp; Hillary. Love it @patrickhealynyt https://t.co/Rvq73ChPSM
DanielAPfister|nytimes|0.8519|0.0|0.491|0.509|Great feature on Madonna &amp; Hillary. Love it @patrickhealynyt https://t.co/Rvq73ChPSM
wear_here|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
iservhomes|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
Pamelapilates|_Proud_American|0.0|0.0|1.0|0.0|RT @_Proud_American: WE FOUND IT! The Video George Soros &amp; Hillary Clinton Tried To Bury! - YouTube https://t.co/Iz9WeknVDW
Pamelapilates|youtube|0.0|0.0|1.0|0.0|RT @_Proud_American: WE FOUND IT! The Video George Soros &amp; Hillary Clinton Tried To Bury! - YouTube https://t.co/Iz9WeknVDW
babysgramma|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
luvmom8702|janet_yackle|-0.3612|0.167|0.739|0.094|"RT @janet_yackle: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/MoUSXY0OP6 via @crooksandlia"
luvmom8702|crooksandliars|-0.3612|0.167|0.739|0.094|"RT @janet_yackle: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/MoUSXY0OP6 via @crooksandlia"
JT4Mets4Arsenal|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/GDeHyTXAio via @Change
JT4Mets4Arsenal|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/GDeHyTXAio via @Change
conservtivegurl|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
deejay90192|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
zaproffo|PeterDoljanin1|-0.4588|0.5|0.5|0.0|@PeterDoljanin1 @American1765 Sorry to disappoint you...https://t.co/63F81u5Mla
zaproffo|independent|-0.4588|0.5|0.5|0.0|@PeterDoljanin1 @American1765 Sorry to disappoint you...https://t.co/63F81u5Mla
photo4art|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
photo4art|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
hnvance40|PeakOfTruth|0.25|0.124|0.677|0.199|RT @PeakOfTruth: Anyone who honestly believes Russia is responsible for #Hillary getting rolled is 2 dumb to continue to draw oxygen https:
AndreFrato|An0nKn0wledge|-0.6739|0.171|0.829|0.0|RT @An0nKn0wledge: THERE IS MORE EVIDENCE OF ALIENS EXISTING THEN THE RUSSIANS HACKING THE ELECTION.. BTW THE ELECTION FRAUD SO FAR ALL IN
xavvypls|twitter|-0.7579|0.302|0.698|0.0|Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure w https://t.co/0szFszOdBd
Ny1david|ibtimes|0.0|0.0|1.0|0.0|Hmmm...https://t.co/QvNiASOjFs
MARGARETFlana18|IdiotDems|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
MARGARETFlana18|t|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
SoBlackAndBlue|twitter|0.0|0.0|1.0|0.0|As opposed to the political juggernauts of Hillary and her team. https://t.co/YnTcsHjLsL
ShaftonP|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
BonnieLCollins3|DemocratCespool|-0.4939|0.158|0.842|0.0|RT @DemocratCespool: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #clintonfoundation http
MacMoney|UberFactsNiggas|0.0|0.0|1.0|0.0|RT @UberFactsNiggas: Hillary Clinton and Snoop Dogg now follow each other on Twitter.
KandorKarteh|kylegriffin1|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
KandorKarteh|theatlantic|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
pinkyfloyd1213|MrDane1982|0.1007|0.161|0.714|0.125|"RT @MrDane1982: 40 yrs of fighting for us, this time we fight for her until she have enough ground to stand on! The best thing Hillary can"
Tish47Patricia|hale_razor|-0.1573|0.125|0.772|0.103|RT @hale_razor: Putin is so brilliant he masterminded Hillary getting 3M more votes than Trump but still lose the election by almost 75 ele
Madam_Nyobi|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
himm7|CarlNyberg312|-0.5574|0.247|0.753|0.0|RT @CarlNyberg312: Hillary Democrat narrative:1. Hillary lost due to sexism.2. Bernie would have lost too. https://t.co/1Qg1MVF0S3
himm7|twitter|-0.5574|0.247|0.753|0.0|RT @CarlNyberg312: Hillary Democrat narrative:1. Hillary lost due to sexism.2. Bernie would have lost too. https://t.co/1Qg1MVF0S3
PatHarr64573322|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
tx_blue_dot|Petergrand|-0.3818|0.14|0.86|0.0|RT @Petergrand: The founding fathers foresaw this situation and designed an emergency override switch called the #ElectoralCollegehttps:/
VeroPArtist|bennydiego|0.2382|0.0|0.911|0.089|RT @bennydiego: It's funny how Hillary's private server was such a major issue but President-elect talking to world leaders on his private
OccuWorld|mediaite|-0.5267|0.221|0.779|0.0|Former U.S. Ambassador to Russia: Vladimir Putin Wanted Revenge on Hillary Clinton https://t.co/802q1LAtdP
fedagentmark|Roscali|-0.2023|0.192|0.657|0.152|@Roscali @almac8241951 @Broker617 @Adjustedwell HILLARY'S bitch Chuck Todd was schooled on truthful journalism by P https://t.co/hFzjP9oSVM
fedagentmark|twitter|-0.2023|0.192|0.657|0.152|@Roscali @almac8241951 @Broker617 @Adjustedwell HILLARY'S bitch Chuck Todd was schooled on truthful journalism by P https://t.co/hFzjP9oSVM
AmericanMom2|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
AmericanMom2|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
HeysannaHosanna|memnosoncos|0.0997|0.198|0.546|0.256|"RT @memnosoncos: ""But please never stop believing that fighting for whats right is worth it."" HillaryGrace under pressure."
bobbyward2009|FoxNews|-0.5423|0.269|0.627|0.103|@FoxNews Hillary is the simple reason the Democrats lost. You sent someone to a gun fight with a knife. Popular vote means nothing.
Workers4Trump|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
JessiePow|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
slone|twitter|-0.565|0.233|0.767|0.0|WHO DIDN'T?????????? The list of people who despise Hillary is very long! https://t.co/H3YZOroavx
CiaoBebe|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
CiaoBebe|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
Rachelle_jdh|ih8florida|0.0772|0.0|0.885|0.115|"@ih8florida @SigmaRoman @arcadianathina @REDLEAFY777 @glamourizes Americans want Hillary, even the republicans"
goldcamaro|CdnChange|0.5562|0.0|0.626|0.374|"4,832,000 strong and counting! https://t.co/GEPVHi9C5E via @CdnChange"
goldcamaro|change|0.5562|0.0|0.626|0.374|"4,832,000 strong and counting! https://t.co/GEPVHi9C5E via @CdnChange"
mosfoodographer|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
mosfoodographer|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
twilbib1|Alyssa_Milano|-0.8173|0.349|0.651|0.0|@Alyssa_Milano more bullshit from Alyssa girl don't have a life get over it asshole Hillary is a criminal
janet_yackle|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
DemClintonKaine|AdamParkhomenko|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
DemClintonKaine|nydailynews|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
ggprez|CarmineZozzora|-0.5267|0.175|0.825|0.0|RT @CarmineZozzora: Russia didn't conspire to delegitimize and sabotage @realDonaldTrump's candidacy or his victory over Hillary Clinton.
mikew6161|NateSilver538|0.8982|0.0|0.502|0.498|"@NateSilver538 LOL. If Hillary didn't cheat, Bernie would have been the nominee.  Enjoy your fairyland dreams."
CerulloElaine|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
dj4k4000|PolitixGal|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
dj4k4000|twitter|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
naja_studio|twitter|0.296|0.111|0.721|0.168|"McCain is all about himself. I am confused where's loyalty stand, he may have voted for Hillary. https://t.co/sSSFKyyvGx"
MarkHoenig|KansasCity1980|0.0|0.0|1.0|0.0|@KansasCity1980 @Lofty537 @parisi_v @WalshFreedom https://t.co/dBoAeJhtdB
MarkHoenig|politifact|0.0|0.0|1.0|0.0|@KansasCity1980 @Lofty537 @parisi_v @WalshFreedom https://t.co/dBoAeJhtdB
oonasez|peterdaou|-0.7579|0.283|0.717|0.0|RT @peterdaou: I've disagreed with Hillary on several issues. I've said her campaign made mistakes. But I'll ALWAYS reject the claim she's
65intexas|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
heatherEcoast|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
MyPlace4U|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
WaldeckKaren|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Future_Comedian|gourmetspud|-0.7717|0.3|0.7|0.0|"RT @gourmetspud: ""Hillary lost bc fake news"" seems 100x less plausible than ""Hillary lost because she was Democratic Romney in anger-driven"
rmbrice|brandongroeny|-0.5106|0.13|0.87|0.0|RT @brandongroeny: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
TXsnark7|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
TXsnark7|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
yvetoro|RJGatorEsq|0.636|0.0|0.811|0.189|RT @RJGatorEsq: Congratulations to President-Elect #Trump on being #Time's Person of the Year! I assume Hillary came in second. #A
assssssssroight|righteousaxe|-0.7506|0.362|0.542|0.096|@righteousaxe @Khanoisseur @mrp @Green_Footballs jesus christ you people are incapable admitting your faults. hillary sucked. simple truth
bittopper_com|bittopper|0.0|0.0|1.0|0.0|Hillary Clinton 2007 Presidential Decks 2008 Vote Hillary.. #rt2gain #teamfollowback #followback #f4f https://t.co/9Ud0laXMS7
constantino_sam|pinterest|0.1531|0.172|0.623|0.206|If you are voting for Hillary  - ANTI HILLARY POLITICAL BUMPER FUNNY STICKER https://t.co/iMfTmpZKmE
PheroNike|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: #PodestaEmails more proof of Hillary's Russian Connections. ""Grassley Letter"" to Loretta Lynch. #CorruptMedia let this stor"
smell3roses|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
westinghouse565|TrinityNYC|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
westinghouse565|t|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
CerulloElaine|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
saminhim|paulbenedict7|-0.7906|0.333|0.667|0.0|RT @paulbenedict7: #Obamastan's FBI: no need to prosecute Hillary's uranium deal; Obamastan's CIA: Putin is a #Trump lobbyist. Worse than #
TXhistorylover|HillaryClinton|-0.1179|0.209|0.6|0.191|so .@HillaryClinton says the Russians rigged the election for Trump to win. Why? Why would they want Hillary to lose?
ZKondos|ABCPolitics|-0.5423|0.189|0.811|0.0|@ABCPolitics Bipartisan my ass. McCain and Graham the two pawns of the #illuminati and Hillary/Obama surrogates...
roqchrisy|WayneDupreeShow|0.0|0.0|1.0|0.0|"RT @WayneDupreeShow: When Obama spoke with Russia in 2012, he said he would have leverage on hot mic, Hillary hit reset button with Putin.."
PatHarr64573322|nytimes|0.3182|0.0|0.874|0.126|RT @nytimes: How a speech by Madonna about sexism put Hillary Clinton's candidacy in fresh perspective https://t.co/CqLswtts4u https://t.co
PatHarr64573322|nytimes|0.3182|0.0|0.874|0.126|RT @nytimes: How a speech by Madonna about sexism put Hillary Clinton's candidacy in fresh perspective https://t.co/CqLswtts4u https://t.co
syl_pac|Change|0.0|0.0|1.0|0.0|Barack Obama: Make Hillary Clinton A Recess Appointment to SCOTUS - Sign the Petition! https://t.co/9K2ug8BgV8 via @Change
syl_pac|change|0.0|0.0|1.0|0.0|Barack Obama: Make Hillary Clinton A Recess Appointment to SCOTUS - Sign the Petition! https://t.co/9K2ug8BgV8 via @Change
HillaryWasRight|Ifitsthisname|-0.8885|0.418|0.509|0.073|@Ifitsthisname @ValeriaPugliesi @JustEric Kennedy and Hatch both created Hillary. You're version is bullshit and you're an evil liar
bzazzie|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
mariebayarea4|VABVOX|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
mariebayarea4|t|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
SilentDogoode|insider|-0.7717|0.456|0.544|0.0|Conway Getting Death Threats Based on 'Incendiary' Anti-Trump Rhetoric https://t.co/GOltPNJOhJ
GarrigaMelissa|DougHenwood|-0.4588|0.2|0.8|0.0|"@DougHenwood @johnphotos he prob means that Hillary, CIA et all are being hypocritical."
aschops|MarkDiStef|0.0|0.106|0.787|0.106|@MarkDiStef @thomas_violence Odd how he's sure of that when polls started to sour on HRC before Comey came along.https://t.co/gwEAa3VVtR
yg_bates|T_Clark8|0.6077|0.073|0.713|0.214|@T_Clark8 how don't I serve the country. I don't see you giving up all your freedoms so everyone else can have theres. you hillary lover
bfm4440|MMFlint|-0.6966|0.2|0.8|0.0|RT @MMFlint: Have you heard a ONE Dem leader scream about this? Imagine if Cuba hacked in to throw the election to Hillary? What would Repu
RickySi16087724|WEdwarda|-0.5848|0.24|0.76|0.0|RT @WEdwarda: @1stcitizen Kills me that Obama campaigned for Hillary on our dime!
Tymeeks98|mitchellvii|0.4019|0.0|0.847|0.153|"@mitchellvii @JohnFromCranber Didn't Mexico try to help Hillary, by having Mexican citizens infiltrate US election process? "
textifyer59|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: I repeat: I laid out what was going on with Russian campaign, based on leaks from European intel, before election: http"
TRESWORLD|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
nana5greatgrand|American1765|-0.5859|0.231|0.769|0.0|RT @American1765: #SundayMorning Reince Priebus #ThisWeek #FakeNewsRussians didn't tell Hillary Clinton 2 ignore MI &amp; WI. Hillary lost bc
shogunofsin|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
faithbasedplans|CebuSalute|0.5093|0.1|0.687|0.213|RT @CebuSalute: haha! Didn't take long for this SJW &amp; Hillary supporting pin-head to block me. Part of the open-minded journalist crowd. ht
travelanita|FoxNews|0.5574|0.113|0.602|0.286|@FoxNews Why would Russia want to defeat their friend Hillary who sold them US Uranium and is friends with Putin?
olivefotini|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
JMCFRAVA|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
millennialviews|madonna|0.296|0.169|0.584|0.247|"Wow, @madonna upset about being called what she really is. https://t.co/BjdNSwdJDT"
millennialviews|mobile|0.296|0.169|0.584|0.247|"Wow, @madonna upset about being called what she really is. https://t.co/BjdNSwdJDT"
TeresaHutson1|DustinGiebel|-0.4019|0.172|0.828|0.0|RT @DustinGiebel: Hillary hacked the DNC because Trump was hogging all the attention.  #BoltonFalseFlagExcuses
PheroNike|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Jakekerrigan17|NoHoesGeorge|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
Jakekerrigan17|twitter|0.6166|0.0|0.748|0.252|RT @NoHoesGeorge: NEVER MAKE FUN OF HILLARY CLINTON IN FRONT OF FEMALES https://t.co/VvtB0z3L0G
roqchrisy|jimlibertarian|0.4939|0.0|0.856|0.144|"RT @jimlibertarian: Donald Trump only works 4 we the people and America,Hillary Clinton on the other hand is a Chinese/Russian agent,she so"
inglamwetrust|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
CerulloElaine|Lrihendry|-0.4767|0.153|0.764|0.083|"RT @Lrihendry: Folks, we need to get on our knees and thank the Lord for sparing us from the impending socialist hell Hillary would've perp"
3Panda3|HeyTammyBruce|0.4404|0.0|0.861|0.139|"RT @HeyTammyBruce: Of course. We've been dealing w ""secret"" CIA report revealed to a Hillary supporting blog (WaPost) by anonymous sources."
farmgurl3|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
AmericanMom2|RepStevenSmith|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
AmericanMom2|dailycaller|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
BillBillmorris|Old_Bern_Kenobi|-0.7579|0.255|0.745|0.0|RT @Old_Bern_Kenobi: This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of fac
theocintric|TheSantaParty|-0.4939|0.167|0.833|0.0|RT @TheSantaParty: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - https://t.co/jALmHrnlkL
theocintric|vivaliberty|-0.4939|0.167|0.833|0.0|RT @TheSantaParty: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - https://t.co/jALmHrnlkL
Kmich718|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
wendydcoe|ali|-0.4404|0.112|0.888|0.0|RT @ali: The media won't point to a single thing Hillary Clinton believes or has done outside of the email scandal that Americans may have
Kevin_thefuture|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
Kevin_thefuture|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
TheJonFerns|guntrust|0.0|0.0|1.0|0.0|RT @guntrust: Wikileaks: Dana Loesch - Hillary's Middle Eastern Firearms Deals Sent Cash to Clinton https://t.co/QVYT2lZhGR #tcot #ccot #2A
TheJonFerns|lawnews|0.0|0.0|1.0|0.0|RT @guntrust: Wikileaks: Dana Loesch - Hillary's Middle Eastern Firearms Deals Sent Cash to Clinton https://t.co/QVYT2lZhGR #tcot #ccot #2A
Politacs7|twitter|0.0|0.0|1.0|0.0|"Ah, so that's what those UFOs have been doing? Wondered about that. Hillary must be one of them. https://t.co/Ln1VtQ3HUG"
hwholcomb|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
ekite56|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
ekite56|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
wendirogersTV|jonleeanderson|0.6808|0.145|0.578|0.277|RT @jonleeanderson: So the CIA says Kremlin hacked Hillary &amp; leaked intel to help Trump.He won &amp; will name a Putin friend Sec of State. Hav
VFL2013|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
VFL2013|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
garki50|VeBo1991|0.5574|0.07|0.696|0.234|RT @VeBo1991: #Hillary loves #Russia when it's funneling $ into her coffers @SteveBo22 https://t.co/wLVDxZVhu6
garki50|twitter|0.5574|0.07|0.696|0.234|RT @VeBo1991: #Hillary loves #Russia when it's funneling $ into her coffers @SteveBo22 https://t.co/wLVDxZVhu6
andsandoval|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Pennie_Bennie|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
Pennie_Bennie|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
PatHarr64573322|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
PatHarr64573322|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
Ikipr|whalefishery|-0.4019|0.213|0.787|0.0|RT @whalefishery: remember when the russians hacked hillary's motor cortex? https://t.co/Mpaek1vD5n
Ikipr|twitter|-0.4019|0.213|0.787|0.0|RT @whalefishery: remember when the russians hacked hillary's motor cortex? https://t.co/Mpaek1vD5n
fool4thetruth|twitter|-0.717|0.23|0.77|0.0|Hillary is the one tied to Russia!!Why are we even wasting time talking about nonsense that Trump had ties to Russ https://t.co/Iim8WHlv9y
beulahcrusoe|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
ggbootsrock|PolitixGal|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
ggbootsrock|twitter|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
KateGriswold1|movietvtechgeek|0.0|0.0|1.0|0.0|RT @movietvtechgeek: the Hillary Clinton Michael Jackson #FakeNews connection #DonaldTrump #MovieTVTechGeeks https://t.co/fB3dJR9Jsw via @m
KateGriswold1|movietvtechgeeks|0.0|0.0|1.0|0.0|RT @movietvtechgeek: the Hillary Clinton Michael Jackson #FakeNews connection #DonaldTrump #MovieTVTechGeeks https://t.co/fB3dJR9Jsw via @m
JessicaRN1995|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
JessicaRN1995|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
LatinoLa2|BigBobGardner|-0.2373|0.148|0.702|0.15|@BigBobGardner @nytimes I tweeted Trump if you want to check... to bet her and do not cry later... Voter fraud for Hillary
oldschoolvet74|DaysOfTrump|-0.5994|0.196|0.804|0.0|"RT @DaysOfTrump: #AmericaFirst Patriots inside USgov are waging a civil war w international socialists (Hillary, Soros..) that have infiltr"
MariuAntonini|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Oldyella49|WalshFreedom|0.5859|0.0|0.84|0.16|"RT @WalshFreedom: If there was evidence that the Russians helped Hillary win, my fellow conservatives would be yelling for an investigation"
lrnewton1|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
marymac169|PrayerChain4HRC|0.4926|0.0|0.834|0.166|RT @PrayerChain4HRC: People putting their Hillary signs back in their yards-now that's truly claiming the victory! @POTUS
HeysannaHosanna|heatherpeno|-0.5423|0.241|0.759|0.0|RT @heatherpeno: When did Hillary &amp; Bernie make Russia the enemy? https://t.co/RatZnIjcAO
HeysannaHosanna|twitter|-0.5423|0.241|0.759|0.0|RT @heatherpeno: When did Hillary &amp; Bernie make Russia the enemy? https://t.co/RatZnIjcAO
JillybeanButtle|eboldy|-0.2263|0.213|0.787|0.0|RT @eboldy: And this.Do. Not. Forget. This.https://t.co/KeEtGhihQh https://t.co/5mIZjaaRzw
JillybeanButtle|twitter|-0.2263|0.213|0.787|0.0|RT @eboldy: And this.Do. Not. Forget. This.https://t.co/KeEtGhihQh https://t.co/5mIZjaaRzw
allofusfortrump|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
LeenaNevaTuuli|France4Hillary|-0.4003|0.306|0.552|0.141|"@France4Hillary @wtfnewsamerica @CIA Charged with treason + Hillary POTUS + EC voting Hillary, please!"
adiazpi|NewsRepublicans|0.0|0.0|1.0|0.0|". @NewsRepublicans @EjHirschberger Obama fue en los hechos el jefe de campaa de Hillary, y perdi; su imprudencia lo est perdiendo hoy"
TatianaBru|CronkiteSays|-0.3818|0.205|0.697|0.098|RT @CronkiteSays: REAL NEWSWe've completed an extensive analysis into why Hillary lost and have determined Hillary caused Hillary to lose
ChristineDBaker|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
heskipto|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
M_IQ_1|VABVOX|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
M_IQ_1|t|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
Lynda_Montgo|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
donnalburnell|JSavoly|-0.7378|0.308|0.692|0.0|RT @JSavoly: Silvers Election Autopsy And Reason For Hillarys Loss Will INFURIATE Everyone #StollenElection #ComradeTrump  https://t.co/v
donnalburnell|abhinavvadrevu|-0.7378|0.308|0.692|0.0|RT @JSavoly: Silvers Election Autopsy And Reason For Hillarys Loss Will INFURIATE Everyone #StollenElection #ComradeTrump  https://t.co/v
Itsgamedayy|AmericanMex067|0.34|0.093|0.701|0.206|"RT @AmericanMex067: .@jmpalmieri says victory came from giving white supremacists a platform. They endorsed Hillary, not Trump. They still"
infidel_murdoc|twitter|0.0|0.0|1.0|0.0|the biggest contributor to his campaign was the american people. but for hillary was the saudi govt https://t.co/sHoPjbhCQu
truthaddict76|DrTomMartinPhD|0.471|0.13|0.663|0.206|"RT @DrTomMartinPhD: HILLARY WON! Current Lead: 2,835,000 Votes. (tiny little side note: DONALD TRUMP IS GUILTY OF TREASON!!!!).  #AMJoy htt"
Lyzvon|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Len51220995|twitter|0.0|0.0|1.0|0.0|"Then don't put your opinion out there OR ..  Hillary is it you ? What,  Bill left again for #PedoFiles island or o https://t.co/1CzS5lDIu4"
coolcatcris|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Greenologue|ElvisNixon7|0.0|0.0|1.0|0.0|@ElvisNixon7 https://t.co/1ZZrPQw9tR
Greenologue|snopes|0.0|0.0|1.0|0.0|@ElvisNixon7 https://t.co/1ZZrPQw9tR
tietude|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: People weren't concerned about Russia when Hillary was selling them US uranium.#MAGA
fritosandmambas|DeplorableTrain|0.5859|0.0|0.858|0.142|RT @DeplorableTrain: Is it possible that Putin wanted Trump to win because he wanted to keep Russia out of WW3 (which would have happened i
DrewSwa|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
Worldofcraze|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
Worldofcraze|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
Goodnightma|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
PaulaChertok|twitter|0.2263|0.105|0.753|0.142|"You're too kind, Tom. They'd skip the witch trials this time and just burn Hillary at the stake. #Kleptocracy https://t.co/eLjbRY5oPS"
amrightnow|twitter|0.0|0.0|1.0|0.0|Hillary Clinton should be in Jail Not on the campaign Trail #realdonaldtrump #military #army #navy #usmc https://t.co/wxjXy80muy
jetsxoxo|Iam_Canadian|-0.5423|0.251|0.664|0.085|"""Hillary=criminal""- @Iam_Canadian agrees her Saudi endorsements should be prosecuted, Russia is a scapegoat &amp; Palestine is under genoside"
KPanderson|AdamParkhomenko|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
KPanderson|nydailynews|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
LiberalsareIcky|YouTube|0.0|0.0|1.0|0.0|Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!  https://t.co/MywrELyiSI via @YouTube
LiberalsareIcky|youtube|0.0|0.0|1.0|0.0|Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!  https://t.co/MywrELyiSI via @YouTube
nana5greatgrand|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
nana5greatgrand||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
PalinInspiresMe|SarahPalinUSA|-0.631|0.153|0.847|0.0|"RT @SarahPalinUSA: Busted. Obama and Hillary voted ""yes"" on building the wall but attack us for that mission today. Does it do any... https"
shoahnuffin1|JeremyHimli|-0.6369|0.346|0.472|0.181|"@JeremyHimli no, idiot like you think that. That's why you helped Hillary. Makes sense. God you're dumb"
Evertonius|neontaster|0.4215|0.0|0.843|0.157|@neontaster @TonyRoller1 I can't believe Russian hackers railroaded @donnabrazile into sharing @CNN debate questions with Hillary #fakenews
mariecasey1|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: Think bout this: Allied intel servives investigating prez-elect 2 learn if he's Putin stooge in place 2 shatter NATO ht
HillaryWasRight|BresPolitico|-0.5754|0.264|0.627|0.109|"@BresPolitico Only stunning this is entire media isnt calling on electors to pick Hillary, reject this dangerous administration"
wendydcoe|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
frodo3245|asamjulian|-0.6159|0.285|0.611|0.104|RT @asamjulian: Funny watching libs cry about Russian interference (w/ no evidence) that didnt care at all about Hillarys MANY foreign i
Goodnightma|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
KateAnn007|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
dwulke|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
KimbaGross|greenhousenyt|0.0|0.0|1.0|0.0|@greenhousenyt @danspence2006 really but investigating HILLARY 24/7 was what??? BI-partisan?
chris_dziuban|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
chris_dziuban|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
iamdansim|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
ChristophSouza|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
TecReview|tecreview|0.0|0.0|1.0|0.0|As fue como Donald Trump pudo superar a Hillary Clinton en los ltimos das de campaa en Estados Unidos https://t.co/7dgPZzDzhh
noelcbickford|JimmyBear2|-0.3818|0.194|0.806|0.0|"RT @JimmyBear2: Hillary Tried To Warn Us About Russia, But Men On Debate Stage Interrupted (VIDEO) - https://t.co/C1qbCUg6i8"
noelcbickford|occupydemocrats|-0.3818|0.194|0.806|0.0|"RT @JimmyBear2: Hillary Tried To Warn Us About Russia, But Men On Debate Stage Interrupted (VIDEO) - https://t.co/C1qbCUg6i8"
cisco_polo711|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
ajitdatta|charliekirk11|-0.5106|0.13|0.87|0.0|RT @charliekirk11: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
HillDamon2015|patriotsphere|0.0|0.0|1.0|0.0|#Fp2017 #Pic #Afd2017 #Petry2017 #Afd #Pictures #Alternativefurdeutschland #Fraukepetry2017 #Fraukepetry #Frauke20 https://t.co/zwTWouEfcN
IndeCardio|1alice4trump|0.3612|0.0|0.872|0.128|RT @1alice4trump: @davidf4444 @riki7s @vivelafra @ChristiChat  leakd email..hillary wanted to make an example of seth .podestra agree. i im
Zelidasquare|fain_2|0.0|0.0|1.0|0.0|"RT @fain_2: @mitchellvii In the words of corrupt crooked Hillary, At this point what difference does it make!"
tanto_dull|MrTriggles|0.0|0.0|1.0|0.0|RT @MrTriggles: @Hypnogogic_Monk @FailureHatesYou @UAsTopSecret @Lonewolf031 @PatriarchyBear @whitesithmale @Sugar_Tits_Bear @JacobRGuillor
JagbusAnne|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: Think bout this: Allied intel servives investigating prez-elect 2 learn if he's Putin stooge in place 2 shatter NATO ht
JosieNano|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
democracydiva|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
democracydiva||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
MaRicky8675309|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
1isten_up|Vote_American|0.0|0.0|1.0|0.0|RT @Vote_American: Maybe there was Russian intervention. But why weren't Dems so intent on finding out whether Hillary's Private Server was
di8285502|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
dblittlefield|twitter|0.6997|0.0|0.766|0.234|"Oh yeah, and I suppose Hillary ran the cleanest, most honest campaign in history.  Such BS.  You could have run, Jo https://t.co/wIiuM0hD7v"
MatthewHrenak|Forbes|-0.6476|0.306|0.694|0.0|@Forbes and they rallied for Hillary and they loss. See! They are the problem
glennasonly|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
galextaft|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
AmericanMom2|tteegar|-0.5242|0.232|0.67|0.098|RT @tteegar: BREAKING #RussianHackers made Hillary screech like an old crabby grandma &amp; lose the election!Nobody should be fooled! #Fak
DanLMcCaughan|Harry1T6|0.0772|0.11|0.769|0.121|RT @Harry1T6: Impressive how Russian hackers forced Hillary Clinton to say she would put coal miners out of business and raise their taxes.
StoneColdChik|StoneColdChik|-0.5816|0.274|0.726|0.0|RT @StoneColdChik: https://t.co/AVW0Tw5fal guess hill stein is really upset with hillary!!!
StoneColdChik|redstatewatcher|-0.5816|0.274|0.726|0.0|RT @StoneColdChik: https://t.co/AVW0Tw5fal guess hill stein is really upset with hillary!!!
TexMexDesi|Remroum|-0.6597|0.252|0.748|0.0|"RT @Remroum: Hillary Clinton lost the election because she is terrible at life, not because a foreign nation intervened."
PraicD|kylegriffin1|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
PraicD|theatlantic|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
robotbum|reason|-0.765|0.28|0.72|0.0|Hillary Clintons Call for Congress to Do Something About Fake News Epidemic Is a Reminder of How Bad Her... https://t.co/ODVEma61d8
Michelem1998|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
ConservativLuke|unsavoryagents|-0.7019|0.243|0.757|0.0|"RT @unsavoryagents: FOR THE RECORD:I AINT ON THE TRUMP TRAIN! I'M ON THE ""FUCK HILLARY"" CABOOSE!"
snowstorm1944|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
FourCM|jonleeanderson|0.6808|0.145|0.578|0.277|RT @jonleeanderson: So the CIA says Kremlin hacked Hillary &amp; leaked intel to help Trump.He won &amp; will name a Putin friend Sec of State. Hav
TheSantaParty|vivaliberty|-0.4939|0.186|0.814|0.0|Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - https://t.co/jALmHrnlkL
raeohkayy|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
YouKeepTheChang|vnuek|-0.1027|0.111|0.796|0.093|"RT @vnuek: Hillary Clinton is well known con artist. 3 weeks after concession she initiates ""recount""... During Dem primaries, she rigged"
RonCentrelloJr|DailyCaller|0.0|0.0|1.0|0.0|@DailyCaller Obama just getting practice for Hillary...
ActionTime|ActionTime|0.0516|0.162|0.669|0.169|RT @ActionTime: Trump Backs Off Campaign Promises Again &amp; Again:Trump Admits His Threat to Lock Up Hillary Was Total Lie #Resist #RT https:
7tips1|tteegar|-0.5242|0.232|0.67|0.098|RT @tteegar: BREAKING #RussianHackers made Hillary screech like an old crabby grandma &amp; lose the election!Nobody should be fooled! #Fak
CherokeeLair|newsweek|0.0|0.0|1.0|0.0|This is happening~ #NuclearWinterIsComing https://t.co/Hyn1TCwvhw
etara44|JudicialWatch|0.0|0.0|1.0|0.0|RT @JudicialWatch: In this country our leaders are bound by the rule of law. Hillary Clinton must be held accountable for her actions.http
MsPGraceMiles|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
kimberlymontse1|HeyTammyBruce|0.4404|0.0|0.861|0.139|"RT @HeyTammyBruce: Of course. We've been dealing w ""secret"" CIA report revealed to a Hillary supporting blog (WaPost) by anonymous sources."
farmgurl3|brandongroeny|-0.5106|0.13|0.87|0.0|RT @brandongroeny: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
TheWomensWatch|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
PalinInspiresMe|SarahPalinUSA|0.0258|0.118|0.759|0.122|RT @SarahPalinUSA: Liberal young'uns... duped again. Hope their parents aren't shelling out big bucks for an education resulting in... http
Diannarinratmom|WhyOpinion|0.25|0.074|0.795|0.131|RT @WhyOpinion: @MissLizzyNJ WikiLeaks email exposed Hillary's oil pipeline with Qatar &amp; truth about Russia https://t.co/GZ87nbsObQ
Diannarinratmom|twitter|0.25|0.074|0.795|0.131|RT @WhyOpinion: @MissLizzyNJ WikiLeaks email exposed Hillary's oil pipeline with Qatar &amp; truth about Russia https://t.co/GZ87nbsObQ
StoneColdChik|redstatewatcher|-0.5816|0.32|0.68|0.0|https://t.co/AVW0Tw5fal guess hill stein is really upset with hillary!!!
halfdollar54|YouTube|0.0|0.0|1.0|0.0|TRUMP ALL-STAR CONWAY JUST RIPPED HILLARY CLINTON A NEW ONE WITH EPIC RA... https://t.co/kFnDPCgUoI via @YouTube
halfdollar54|youtube|0.0|0.0|1.0|0.0|TRUMP ALL-STAR CONWAY JUST RIPPED HILLARY CLINTON A NEW ONE WITH EPIC RA... https://t.co/kFnDPCgUoI via @YouTube
Millenniumistic|MadameWoo69|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
Millenniumistic|change|0.0|0.0|1.0|0.0|RT @MadameWoo69: Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/TTrq3BfMmc via @Change
Debbie1228Hart1|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
boydmyers|PalmettoMoon214|0.4515|0.113|0.646|0.241|RT @PalmettoMoon214: #ITriedHardBut I can't stop laughing at this clip of Hillary prematurely thinking she won the election.  https://t.co
boydmyers|t|0.4515|0.113|0.646|0.241|RT @PalmettoMoon214: #ITriedHardBut I can't stop laughing at this clip of Hillary prematurely thinking she won the election.  https://t.co
cahulaan|rbaker65708|-0.8482|0.281|0.719|0.0|"@rbaker65708 @Pink22Karen @thinkprogress I am so sick of this shit, why put up with it? What can we do besides petitions etc? Com'on Hillary"
Col_Connaughton|youtube|0.3182|0.0|0.859|0.141|"Truth vs. NEW$, Inc. Sept 15 2016, Fetzer, Bennett, Part 2 https://t.co/rMC9NnpBqU #hillary #clinton #double #911"
flyer74|flyer74|-0.8429|0.335|0.665|0.0|RT @flyer74: MR. FAKE NEWS HIMSELF..........ON THE HILLARY CLINTON FOUNDATION DIVISION OF THE CLINTON CRIME FAMILY PAYROLL....... https://t
flyer74||-0.8429|0.335|0.665|0.0|RT @flyer74: MR. FAKE NEWS HIMSELF..........ON THE HILLARY CLINTON FOUNDATION DIVISION OF THE CLINTON CRIME FAMILY PAYROLL....... https://t
SEH101184|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
rzitka|aquawilki|-0.5096|0.3|0.7|0.0|@aquawilki @CliftonsNotes didn't he promise to jail Hillary.  Now he isn't. Lol.
roqchrisy|DebAlwaystrump|0.5405|0.0|0.776|0.224|RT @DebAlwaystrump: HILLARY SELLS 20% OF USA URANIUM TO RUSSIAWHYDems must not be too worried about Russia sure Russia would want more
sassysassyred|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
gamecocksSecE|heyjoshhaines|-0.8813|0.295|0.705|0.0|".@heyjoshhaines but the info has been leaked and has shown corruotion &amp; collusion by MSM, Hillary,DNC, etc that is very much so wrong doing!"
VegasVictory|vivaliberty|-0.4939|0.176|0.824|0.0|Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.co/3RRDKJkVjy
Kaffe_Takk|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
trickytweeter|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
Chicken_Legz69|YouTube|0.6809|0.0|0.753|0.247|OMG!!!! HILLARY VS TRUMP PRESIDENTIAL DEBATE 10 SUBSCRIBER SPECIAL 50TH VIDEO SPECIAL!!!!!!: https://t.co/4S7AYWzAJq via @YouTube
Chicken_Legz69|youtube|0.6809|0.0|0.753|0.247|OMG!!!! HILLARY VS TRUMP PRESIDENTIAL DEBATE 10 SUBSCRIBER SPECIAL 50TH VIDEO SPECIAL!!!!!!: https://t.co/4S7AYWzAJq via @YouTube
CindyLeinwand12|linkis|0.7184|0.0|0.75|0.25|"In a world where the president makes fun of handicapped people and fat people, how do we proceed with dignity? https://t.co/RvtFKzmz6l"
VivianLeeDavis1|JustNWashington|-0.6166|0.155|0.845|0.0|"@JustNWashington @thehill Doesn't have to mention Hillary, bc Dumbo is a PATHOLOGICAL LIAR &amp; you can take that to the BANK u people will see"
1isten_up|Vote_American|0.0|0.0|1.0|0.0|"RT @Vote_American: @Vote_American If WikiLeaks got to Hillary's Email Private Server, So Did the Russians, China, N Koria, and all others!"
StormSpinning|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
jtinfo|irishspy|0.2732|0.0|0.588|0.412|@irishspy @sistertoldjah Hillary supporter.
winstar1k|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
winstar1k|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
StuNeff|TerriGreenUSA|-0.3612|0.111|0.889|0.0|"RT @TerriGreenUSA: Hillary was careless with her many cell phones and emails. And this happened under Obama's watch, not under a Republican"
MikeTruck62|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
DonnaDeCicco1|Dr_of_Nursing|0.6124|0.0|0.762|0.238|"RT @Dr_of_Nursing: #Treason disqualifies #Trump from being PEOTUS, #ElectoralCollege can easily resolve the issue by choosing #Hillary http"
SiberiaCat3|BrianWestrate|-0.4939|0.168|0.769|0.063|.@BrianWestrate @denadecamp Pls don't vote for Trump. He will destroy the GOP. Hillary works with ALL. #FlipThe37 https://t.co/hGntPGhuox
SiberiaCat3|chicagotribune|-0.4939|0.168|0.769|0.063|.@BrianWestrate @denadecamp Pls don't vote for Trump. He will destroy the GOP. Hillary works with ALL. #FlipThe37 https://t.co/hGntPGhuox
MyPlace4U|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
MyPlace4U|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
theerinmaher|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
CerulloElaine|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
benitah_summers|Rabiddogg|0.4404|0.0|0.879|0.121|RT @Rabiddogg: @SheriffClarke @realDonaldTrump is it safe to assume Hillary can see her own reflection if she stands in front of a mirror?
foothands|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
MicheleWeiss69|TrumpSuperPAC|-0.5423|0.137|0.863|0.0|"RT @TrumpSuperPAC: If Russia is the enemy, why isn't anyone looking into why #Hillary sold 20% of our American Uranium to Russia? #SecretCI"
StillBernin|ojoscriollos|-0.8269|0.421|0.418|0.161|RT @ojoscriollos: Isn't it great when Hillary supporters &amp; someone they've derided as dangerous RWNJ agree are allies in a propaganda war a
hnvance40|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
kwknox50|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/1gh1HI1kL4
MCGA2019|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
Old_Bern_Kenobi|twitter|-0.7579|0.277|0.723|0.0|This is how far Hillary's sycophants have sunk: Blaming fast food workers for Hillary's failure without a shred of https://t.co/7gTWGx9mQx
tgranillo|WalshFreedom|0.5859|0.0|0.84|0.16|"RT @WalshFreedom: If there was evidence that the Russians helped Hillary win, my fellow conservatives would be yelling for an investigation"
TroyCoby|TroyCoby|-0.6705|0.244|0.756|0.0|RT @TroyCoby: Hillary Clinton has lost mostly because she is what she is - the arrogant limo liberal elite... https://t.co/PFpR3DQeTD
TroyCoby|twitter|-0.6705|0.244|0.756|0.0|RT @TroyCoby: Hillary Clinton has lost mostly because she is what she is - the arrogant limo liberal elite... https://t.co/PFpR3DQeTD
SEH101184|emzorbit|-0.4215|0.128|0.872|0.0|RT @emzorbit: @ezlusztig @CNNPolitics And somebody needs to get that crooked toothed Giuliani in a chair and under freaking oath. https://t
SEH101184||-0.4215|0.128|0.872|0.0|RT @emzorbit: @ezlusztig @CNNPolitics And somebody needs to get that crooked toothed Giuliani in a chair and under freaking oath. https://t
LyleELong|DineshDSouza|-0.7579|0.365|0.539|0.095|RT @DineshDSouza: .@HillarysAmerica revealed the truth about Hillary and helped avert disaster. Commemorate her historic defeat: https://t.
LyleELong||-0.7579|0.365|0.539|0.095|RT @DineshDSouza: .@HillarysAmerica revealed the truth about Hillary and helped avert disaster. Commemorate her historic defeat: https://t.
Worldofcraze|Change#|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/HIdztiSuIQ via @Change#
Worldofcraze|linkis|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/HIdztiSuIQ via @Change#
bluebonnetbunny|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
TereseForstbau1|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
JeffersonsNotes|westernlvr|-0.3818|0.212|0.68|0.108|"@westernlvr @WalshFreedom No, they were gross. But a) they were legitimately charitable, and b) Hillary wasn't president. Focus on now?"
hwymanric10|Str8Grandmother|-0.7269|0.289|0.711|0.0|RT @Str8Grandmother: Former US Ambassador: Russia Hacked The Election To Get Revenge Against Hillary Clinton [VIDEO] https://t.co/SOE1agr9XO
hwymanric10|joemygod|-0.7269|0.289|0.711|0.0|RT @Str8Grandmother: Former US Ambassador: Russia Hacked The Election To Get Revenge Against Hillary Clinton [VIDEO] https://t.co/SOE1agr9XO
AleciaWarrenXO|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
PalinInspiresMe|SarahPalinUSA|0.0|0.0|1.0|0.0|RT @SarahPalinUSA: Rush reminds us ---&gt; https://t.co/VdGq41JjmZ https://t.co/BV9NwoEYvq
PalinInspiresMe|youngcons|0.0|0.0|1.0|0.0|RT @SarahPalinUSA: Rush reminds us ---&gt; https://t.co/VdGq41JjmZ https://t.co/BV9NwoEYvq
suzykq5|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
John132941831|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
Magilla7|DaysOfTrump|-0.5994|0.196|0.804|0.0|"RT @DaysOfTrump: #AmericaFirst Patriots inside USgov are waging a civil war w international socialists (Hillary, Soros..) that have infiltr"
johnthepiper|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
melinda118|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
carloshiatt|JBurtonXP|0.6597|0.0|0.779|0.221|"RT @JBurtonXP: If Russia wanted to influence the election, they should've just donated millions to Hillary like all the respectable foreign"
DJT_ChosenbyGod|attentionmustbe|0.0|0.0|1.0|0.0|RT @attentionmustbe: Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!    https://t.co/X81oHLk56F via @YouTube
DJT_ChosenbyGod|youtube|0.0|0.0|1.0|0.0|RT @attentionmustbe: Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!    https://t.co/X81oHLk56F via @YouTube
LatestComPols|latest|-0.6115|0.235|0.765|0.0|Harvard Study: Hillary Clinton Received The Most Negative Coverage in 2016 Campaign https://t.co/CWCAcciZLK https://t.co/29iBjidjYp
shayne571|sullivanamy|0.0|0.0|1.0|0.0|"RT @sullivanamy: That was Joel Benenson's take at U. Chicago a few wks ago. Headlines all scanned as ""emails,"" or ""just more Hillary corrup"
Hotmess_Mello|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
chantellym|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
flyer74|flyer74|0.7885|0.0|0.683|0.317|RT @flyer74: YES IT IS TRUE OBAMA HELPED FORM ISIS ALONG WITH HILLARY CLINTON......GOOD GOING IDIOTS... https://t.co/1ArbKPbg8Z
flyer74|twitter|0.7885|0.0|0.683|0.317|RT @flyer74: YES IT IS TRUE OBAMA HELPED FORM ISIS ALONG WITH HILLARY CLINTON......GOOD GOING IDIOTS... https://t.co/1ArbKPbg8Z
JCCentCom|jtLOL|0.0609|0.082|0.828|0.09|RT @jtLOL: I'll put it like this: Comey wouldn't have needed to send that letter if Hillary Clinton hasn't been so lawless and paranoid. ht
DaeshPussy|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
CocoThePatriot|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
photo4art|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: What if the election hadn't been hacked?What if Hillary hadn't stole the nomination?What if Obama hadn't given rise to
RepublicanPN|twitter|0.126|0.113|0.687|0.199|"You want to know how sick Main Stream Media is just look at this video! Hillary, Obama, only God can forgive you now https://t.co/oyC9cWOOYl"
kldreams61|arian0027|-0.8126|0.355|0.576|0.07|"RT @arian0027: Are you that ignorant, no machines were hacked. Hillary was exposed, and we on Twitter pushed for the truth the lying MSM fa"
kingvideo123|HumanistReport|-0.6705|0.2|0.8|0.0|"RT @HumanistReport: If Hillary Clinton was ever going to denounce fake news, she should have done it after it made her falsely believe Iraq"
perry1949|GrayConnolly|-0.2263|0.136|0.769|0.095|"RT @GrayConnolly: ""Russians forced Hillary to set up Clinton Foundation that accepted Russian money for State Dept favours""...or something"
YosefBorgen|breitbart|-0.508|0.202|0.798|0.0|Holy Cow! ! Report: Hillary Clinton Spent $1.2 Billion to Lose 2016 Election. https://t.co/vROojLaQI5 https://t.co/mk4EBdU4ev
mekmtl|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
AndreFrato|rtyson82|-0.5423|0.304|0.696|0.0|"RT @rtyson82: Hillary still has bad judgment, I see... https://t.co/SK6YONjN7y"
AndreFrato|twitter|-0.5423|0.304|0.696|0.0|"RT @rtyson82: Hillary still has bad judgment, I see... https://t.co/SK6YONjN7y"
loveboat_SANK|twitter|0.0|0.0|1.0|0.0|2 GOP HILLARY CUCKS ! https://t.co/hgzGHBBr8g
Diannarinratmom|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Lisela36Graham|OnlyTruthReign|-0.4574|0.232|0.67|0.098|RT @OnlyTruthReign: @dilemmv @NancyPelosi yep no backbone! Russia Russia Russia gave Hillary $145Mill then #RussiaHackers hacked the electi
SiberiaCat3|candynoble|0.0|0.0|1.0|0.0|.@candynoble We the people have spoken. 2 million more votes for Hillary. #HonorPopularVote #MoralElectors https://t.co/jvinMowiss
SiberiaCat3|twitter|0.0|0.0|1.0|0.0|.@candynoble We the people have spoken. 2 million more votes for Hillary. #HonorPopularVote #MoralElectors https://t.co/jvinMowiss
Syr829|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
OrpheusDescent|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
OrpheusDescent|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
ftabs1931|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
rstantono|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
BelisaDavis|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
zombieninja420|softwarnet|-0.2732|0.091|0.909|0.0|"RT @softwarnet: ""FBI and CIA""Podesta was warned in 2008 to use encryption, Hillary didn't, DNC didn't, Obama's OPM didn't - those who igno"
Valeriegromes16|btrwkart|0.0|0.0|1.0|0.0|@btrwkart @kiddle https://t.co/Kpi03JGKSX
Valeriegromes16|townhall|0.0|0.0|1.0|0.0|@btrwkart @kiddle https://t.co/Kpi03JGKSX
Bane1349|PolitixGal|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
Bane1349|twitter|-0.5147|0.27|0.73|0.0|RT @PolitixGal: This Michigan crowd is WHY HILLARY LOST! https://t.co/mofoGRjQQO
flajeffreyt|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
jsirwin67|original|-0.5994|0.494|0.506|0.0|Hillary is a war monger https://t.co/Id3MZlVOyT
carwizrd|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
johnthepiper|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
1carpediem2016|realjunsonchan|0.4076|0.133|0.632|0.235|"RT @realjunsonchan: -@KellyannePolls completely rekts Rotten Hillary. Lol. This is how America should be governed, spend less, win more. Ni"
elizabethkap|VABVOX|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
elizabethkap|t|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
Psalm11813|redsteeze|0.0|0.0|1.0|0.0|RT @redsteeze: Russia wanted Trump. You know who else wanted Trump? Hillary &amp; our media. All three got what they wanted.
KeelinMadden|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
KeelinMadden|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
Anfoooey|realjunsonchan|0.4076|0.133|0.632|0.235|"RT @realjunsonchan: -@KellyannePolls completely rekts Rotten Hillary. Lol. This is how America should be governed, spend less, win more. Ni"
LauraEmilyPDX|ericgrant|0.0|0.0|1.0|0.0|RT @ericgrant: The takeaway from all this Russian news: everyone should hire the person who set up Hillary's impenetrable email server.
last2brake|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
tdortchlee|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
Andryushallc|JerryT87|0.0|0.0|1.0|0.0|RT @JerryT87: @LeahR77 @AppSame This is what Hillary and gang had planned for us. Bet on it.
WamplerJim|Evan_McMullin|0.5256|0.0|0.825|0.175|@Evan_McMullin @realDonaldTrump a 1000 times more loyal than u and that skank Hillary .. ur 15 minutes are over
GodandtheBear|twitter|-0.7044|0.292|0.708|0.0|What about we don't want Hillary don't you understand? Try all you want you can't make me feel shame for her loss e https://t.co/fAliinPLlJ
clark7950|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: People weren't concerned about Russia when Hillary was selling them US uranium.#MAGA
jwire|bocavista2016|0.0|0.0|1.0|0.0|RT @bocavista2016: Hillary ILLEGALLY sold Russia uranium for NUKESYet Putin/@realDonaldTrump bromance is the Nat Sec threat?https://t.c
jwire||0.0|0.0|1.0|0.0|RT @bocavista2016: Hillary ILLEGALLY sold Russia uranium for NUKESYet Putin/@realDonaldTrump bromance is the Nat Sec threat?https://t.c
theonegenegreen|AtlTeaPartyLove|-0.5267|0.167|0.833|0.0|RT @AtlTeaPartyLove: Hillary Clinton is a danger to everyone rights when she unleash Syrian Rapefugees on our soil https://t.co/CvJBwbjacL
theonegenegreen|twitter|-0.5267|0.167|0.833|0.0|RT @AtlTeaPartyLove: Hillary Clinton is a danger to everyone rights when she unleash Syrian Rapefugees on our soil https://t.co/CvJBwbjacL
writeinussenate|DailyCaller|0.0|0.0|1.0|0.0|@DailyCaller @bzazzie More than hillary and merkel??
1Gadsdenflag2|ed_hooley|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
1Gadsdenflag2|truthfeed|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
ReaganCoalition|fiscalconservatives|0.0|0.0|1.0|0.0|REVEALED  The Hillary Aide Who KNEW It Was All Over https://t.co/pBxUGkdoYl
tonic516|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
oklegacy|pambesteder|0.4404|0.0|0.861|0.139|RT @pambesteder: Didn't Hillary and Obama push the RESET button with Russia because THEY wanted a better relationship with them?
Cc54518746C|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
photo4art|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
annettedufresne|Chemzes|0.0|0.0|1.0|0.0|RT @Chemzes: Me when somebody asks for my thoughts on Hillary Clintonhttps://t.co/VlFIAYCc4K
TrumptheGOP|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
sancusbook|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
curiously_yours|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
jjmikemike|"CNN,"|-0.3182|0.223|0.777|0.0|"Just a reminder from @CNN, from before Hillary lost. https://t.co/xg0c0XllYJ"
jjmikemike|twitter|-0.3182|0.223|0.777|0.0|"Just a reminder from @CNN, from before Hillary lost. https://t.co/xg0c0XllYJ"
debelwar|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
TerriGreenUSA|twitter|-0.3612|0.116|0.884|0.0|"Hillary was careless with her many cell phones and emails. And this happened under Obama's watch, not under a Repub https://t.co/Ok8DxvwVqB"
michelekirkBPR|twitter|-0.4019|0.124|0.876|0.0|"Dem gov. of Virginia recalls omen that spelled doom for Hillary, and it has to do with his chickens https://t.co/5VukS6bAr4"
ScreenCaffeen|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
gscarroll47|Patrici15767099|-0.6908|0.213|0.787|0.0|"RT @Patrici15767099: If Dems big donors are stupid enough to believe Hillary lost the election b/c of Russian influence, they deserve to lo"
rgreen00|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
HillaryBCrooked|LadyPatriot2000|-0.2225|0.161|0.718|0.121|"RT @LadyPatriot2000: Hilarious that these Lefties still aren't over it! Hillary sucked from day 1, still does! https://t.co/kTjTSN9DVQ"
HillaryBCrooked|twitter|-0.2225|0.161|0.718|0.121|"RT @LadyPatriot2000: Hilarious that these Lefties still aren't over it! Hillary sucked from day 1, still does! https://t.co/kTjTSN9DVQ"
TheOneLadyEagle|ReversingASD|-0.25|0.215|0.61|0.175|"RT @ReversingASD: @FoxNews just like Hillary playing the ""Russian card"" &amp; ""fake news card"" to avoid #PayToPlay  indictment @dtrumpnation @"
SiberiaCat3|kyhm1024|0.3818|0.0|0.794|0.206|.@kyhm1024 Take note that Hillary helps children. #FlipThe37 #MoralElectors https://t.co/OxjphTSP7o  https://t.co/Ld8fZcvbuV
SiberiaCat3|gothamist|0.3818|0.0|0.794|0.206|.@kyhm1024 Take note that Hillary helps children. #FlipThe37 #MoralElectors https://t.co/OxjphTSP7o  https://t.co/Ld8fZcvbuV
KerryOtis|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
ZRODWN|YoungDems4Trump|-0.1531|0.082|0.918|0.0|RT @YoungDems4Trump: WikiLeaks Emerges from the Shadows to Expose Stephen Colbert &amp; Hillary's Clinton Global Initiative Ties- @LeahR77 ht
kimberlymontse1|TravisRuger|-0.5994|0.178|0.822|0.0|RT @TravisRuger: Since when did dems start wanting war with Russia so much?   #AMJoy  #imstillwithher #60Minutes #maddow #inners https://t.
kimberlymontse1||-0.5994|0.178|0.822|0.0|RT @TravisRuger: Since when did dems start wanting war with Russia so much?   #AMJoy  #imstillwithher #60Minutes #maddow #inners https://t.
Magilla7|DrMartyFox|0.0|0.0|1.0|0.0|RT @DrMartyFox: We Do Have Evidence Of #RussianMeddlingThe Uranium Deal #Putin Wanted #Hillary To Be President So He Could Make More
poliannesez|CitizensFedUp|0.2023|0.0|0.872|0.128|"RT @CitizensFedUp: Hillary could have legal right to challenge electoral college system and be next US president, says law professor https:"
kierobar|Tis4Ta|-0.1779|0.182|0.657|0.161|"RT @Tis4Ta: Still no lead in Seth Rich death, he work for the government. They should be looking with a fine tooth comb, But for Hillary ev"
LaVerneWright13|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
LaVerneWright13||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
shelbysbroccoli|WalshFreedom|0.5859|0.0|0.84|0.16|"RT @WalshFreedom: If there was evidence that the Russians helped Hillary win, my fellow conservatives would be yelling for an investigation"
imissguinness|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
imissguinness||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
bait51|Tis4Ta|-0.743|0.221|0.708|0.071|"RT @Tis4Ta: I agree with you, &amp; I am mad as hell with why Hillary is not in jail. did she paid everyone off or have deep secrets on them, w"
oklegacy|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
rgreen00|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
rgreen00||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
JulianitaSj|jonleeanderson|0.6808|0.145|0.578|0.277|RT @jonleeanderson: So the CIA says Kremlin hacked Hillary &amp; leaked intel to help Trump.He won &amp; will name a Putin friend Sec of State. Hav
CpturCre8Studio|charliekirk11|-0.5106|0.13|0.87|0.0|RT @charliekirk11: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
ChristophSouza|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
infidel_murdoc|twitter|0.25|0.056|0.847|0.097|your talking about the pay for play when hillary was the SOS. she sold position at a price. it was publish at wikil https://t.co/JLqlvrMAMG
carolinefili|charliekirk11|0.0|0.0|1.0|0.0|"RT @charliekirk11: New evidence shows Russian hackers changed Hillary's speech to include the words ""deplorable and irredeemable"" #FakeNe"
PoliticsToday_|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
kathyschmidt12|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
punkcurmudgeon|Hedge76|-0.765|0.266|0.734|0.0|"RT @Hedge76: Here's the thing: Hillary is crap and she lost a gimme election.  Having said that, we basically elected the Meteor of Doom to"
ChristophSouza|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: The Democrats all debate who's going to get out of Hillary's way first, except for VERMONT'S OWN BERNIE SANDERS, who...get"
TallManShort|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
RealJimPeterson|nia4_trump|-0.7096|0.258|0.742|0.0|RT @nia4_trump: Hillary blames Russia &amp; #FakeNews for her lossReality Check it was the Scandals Corruption Collusion &amp; Divisivenesshttps:
groworx|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
XXXGlassSexToys|change|0.8047|0.0|0.453|0.547|PLEASE SIGN AND RE-TWEET! THANKS EVERYONE! ;-)https://t.co/Cyk9CcAk2d https://t.co/pstowpdZsS
Butch1717|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
gianghoang1705|youtube|0.0|0.0|1.0|0.0|Ti  thch video https://t.co/VFcmeYe1h1 The Second Presidential Debate: Hillary Clinton And Donald Trump (Full Debate) | NBC
News4Newsman|TrumpSuperPAC|-0.7772|0.244|0.756|0.0|RT @TrumpSuperPAC: We came close to the apocalypse with this raving lunatic! #Hillary wants to censor all media! Who's the Nazi now? https:
dawnzer61|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
dawnzer61|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
starlady24|CapitalismCures|0.3612|0.1|0.706|0.193|RT @CapitalismCures: the same people refusing accept Trump as president were yelling that everyone needs to accept the results when they th
rharrisonfries|FrankLuntz|-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
rharrisonfries||-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
typserv|MarthaLivingmar|-0.1134|0.123|0.774|0.103|"RT @MarthaLivingmar: @mitchellvii @DonWeldy And that is because the problems are never their fault, just ask Obama or Hillary."
opelikacreek|gerfingerpoken|0.0772|0.149|0.683|0.168|RT @gerfingerpoken: Did IRS Leak Trump Returns 2 Help Hillary? https://t.co/EWkqWLPAQNAmerican Thinker https://t.co/L7h6rlr1le https://t.
opelikacreek|t|0.0772|0.149|0.683|0.168|RT @gerfingerpoken: Did IRS Leak Trump Returns 2 Help Hillary? https://t.co/EWkqWLPAQNAmerican Thinker https://t.co/L7h6rlr1le https://t.
rgreen00|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
RebeccaKovalich|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
RebeccaKovalich||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
dwulke|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
thalsey51|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
thalsey51||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
HillarysPurse|ComfortablySmug|0.0|0.0|1.0|0.0|"@ComfortablySmug @WalshFreedom Soros (Hillary proxy) meddled with Ukraine elections. Putin was ""Hey"" And we were all ""Whaaa?"""
Sioflynn|Im_ConnorKelley|0.5719|0.0|0.73|0.27|RT @Im_ConnorKelley: @realDonaldTrump @NBCNightlyNews @CNN Hillary won by 2.83 million votes
jsirwin67|original|0.0|0.0|1.0|0.0|https://t.co/Id3MZlVOyT
thickmick59|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
KenMeyer91|mediaite|0.0|0.0|1.0|0.0|Former U.S. Ambassador to Russia: Vladimir Putin Wanted 'Revenge' on Hillary Clinton https://t.co/KO90SKaRuC
mikew6161|DrMartyFox|0.0|0.0|1.0|0.0|RT @DrMartyFox: We Do Have Evidence Of #RussianMeddlingThe Uranium Deal #Putin Wanted #Hillary To Be President So He Could Make More
IBDeb2|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
OriginalVader1|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
OriginalVader1|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
hmrstrm45|SheriffClarke|0.4404|0.0|0.884|0.116|RT @SheriffClarke: This is priceless. I would have paid good money to have been on a conference call hook-up when she made this call. https
cala_1111|truthfeed|-0.5319|0.209|0.791|0.0|This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/zXFrE2Pvg7
GreatNikolajs|Heypag|-0.7003|0.284|0.588|0.127|@Heypag But I think you would rather come up with a lame excuse on how Hillary lost than actually accept that she was a shitty candidate.
linos2015|tonywoody1574|-0.3734|0.217|0.654|0.129|RT @tonywoody1574: @KellyannePolls @nypost it's so funny the left says Russia made Hillary lose Hillary and her EMAILS on her illegal SERVE
tobyonekonobe|MissMandi00|-0.25|0.152|0.738|0.111|"RT @MissMandi00: No.If you're convinced #Hillary is corrupt, flawed, unlikable, &amp; dishonest, you're more in touch w/reality than +/-63 mil"
Freedom1776__|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
Freedom1776__|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
Shalom555222|RepStevenSmith|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
Shalom555222|dailycaller|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
Millenniumistic|1DianeMarie|0.4215|0.11|0.675|0.215|RT @1DianeMarie: @calminsensehypn @DefraudTheVote NO. We Want Hillary Rodham Clinton ONLY. She WON. We deserve to HAVE Her as OUR #MadamePr
dustyfingertips|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
Nan33S|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
teresarc17|ed_hooley|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
teresarc17|truthfeed|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
geoff_deweaver|LoriRMixson|-0.7269|0.319|0.681|0.0|Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/j0iJ78yMVo cc @LoriRMixson @LouDobbs
geoff_deweaver|nytimes|-0.7269|0.319|0.681|0.0|Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/j0iJ78yMVo cc @LoriRMixson @LouDobbs
rm1268|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
RedVote2016|5Against1Eight3|-0.1027|0.195|0.625|0.18|"@5Against1Eight3 God showed them what a baby could understand. If they still choose people like Hillary Clinton, they're lost. Their problem"
RebeccaKovalich|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
NickMarsillo|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
NickMarsillo|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
MyPupVoted|TrumpSuperPAC|-0.4588|0.167|0.833|0.0|"RT @TrumpSuperPAC: The man who hacked #Hillary's personal emails and is currently in prison gave a statement to the legacy media, but they"
Mark_Peabod1|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
Mark_Peabod1|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
ChrisSl66335686|KellyannePolls|-0.5423|0.171|0.829|0.0|@KellyannePolls Hillary didn't have you kicking ass on every talk show and media outlet in the nation https://t.co/ptrcCfGsXh
ChrisSl66335686|twitter|-0.5423|0.171|0.829|0.0|@KellyannePolls Hillary didn't have you kicking ass on every talk show and media outlet in the nation https://t.co/ptrcCfGsXh
mmsahaj|javaguysammckee|0.0|0.0|1.0|0.0|RT @javaguysammckee: @JackPosobiec But they don't mind that Hillary let Putin have control of 20% of world uranium production in exchange f
CherylHodge13|aworldoftruth|-0.2732|0.11|0.89|0.0|RT @aworldoftruth: Hillarys Russian Hack Hoax: The Biggest Lie of This Election Season FBI and CIAhttps://t.co/rIZL9OAKmK via @grtvne
ProChoiceKills|LauraLeeBordas|0.3254|0.151|0.584|0.265|RT @LauraLeeBordas: BOMBSHELL - Journalist Confirms Media Created THIS Fake News Story to HELP Hillary https://t.co/nWt9ERE6Am
ProChoiceKills|angrypatriotmovement|0.3254|0.151|0.584|0.265|RT @LauraLeeBordas: BOMBSHELL - Journalist Confirms Media Created THIS Fake News Story to HELP Hillary https://t.co/nWt9ERE6Am
6353a95c845e426|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
WakeUpCanada1|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
OccupyEnlighten|LAProgressive|0.0|0.0|1.0|0.0|"RT @LAProgressive: Music, Politics, and Hillary https://t.co/wHEldAnzh6 #Feelthebern #Hillaryclinton #Trumptweet https://t.co/GAwxyjUTzw"
OccupyEnlighten|laprogressive|0.0|0.0|1.0|0.0|"RT @LAProgressive: Music, Politics, and Hillary https://t.co/wHEldAnzh6 #Feelthebern #Hillaryclinton #Trumptweet https://t.co/GAwxyjUTzw"
IrishSix1|bad_bad_bernie|-0.1828|0.148|0.738|0.114|RT @bad_bad_bernie: It wasn't the Republicans attacking Hillary that destroyed the Democratic Party.It was the Democrats defending Hillar
Megan_Hafer|Andrew_Hafer|0.3182|0.0|0.566|0.434|"@Andrew_Hafer Calm down, Hillary"
LAangel49|rodneyawilli|-0.4184|0.134|0.866|0.0|RT @rodneyawilli: @kabtlc @TerranomaLead @chuckwoolery Oh the Hypocrisy!!  Imagine if Hillary refused to release her tax returns while Trum
Groughy|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
theo1972|TrumpsDisciple|0.4986|0.112|0.585|0.303|RT @TrumpsDisciple: Thank goodness that Hiterly didn't win. The democrat white supremacist elites baking her would of been chanting Hail Hi
JulieTu52053648|SiessChris|-0.7964|0.336|0.664|0.0|RT @SiessChris: Nope. They were too busy making shit up to cover Hillary's fat ass. https://t.co/OevhAUkfbJ
JulieTu52053648|twitter|-0.7964|0.336|0.664|0.0|RT @SiessChris: Nope. They were too busy making shit up to cover Hillary's fat ass. https://t.co/OevhAUkfbJ
fool4thetruth|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: #PodestaEmails more proof of Hillary's Russian Connections. ""Grassley Letter"" to Loretta Lynch. #CorruptMedia let this stor"
ErickaMinger|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
PeterPeterson95|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
TimBroderick|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
TimBroderick||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
janiceponchak|FreedomChild3|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
janiceponchak|t|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
Stephynb|ParentofSam1|0.0|0.0|1.0|0.0|"RT @ParentofSam1: @USA_First_2016 @kurteichenwald https://t.co/61G4YuKKoT 4,828,260 signatures now... https://t.co/erKnbGPCJ4"
Stephynb|change|0.0|0.0|1.0|0.0|"RT @ParentofSam1: @USA_First_2016 @kurteichenwald https://t.co/61G4YuKKoT 4,828,260 signatures now... https://t.co/erKnbGPCJ4"
PatPatojson|softwarnet|-0.2732|0.091|0.909|0.0|"RT @softwarnet: ""FBI and CIA""Podesta was warned in 2008 to use encryption, Hillary didn't, DNC didn't, Obama's OPM didn't - those who igno"
Joymar27|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
FactsVsOpinion|ReinaA808|-0.2732|0.084|0.916|0.0|RT @ReinaA808: @RadioFreeTom I voted for Hillary cos I knew Trump was going to give Wall St. and the 1% total power. Bernie warned us about
News4Newsman|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
polyglotme|shayne571|-0.4215|0.149|0.851|0.0|@shayne571 @NoyzeSmythe @4everNeverTrump @caliwaterman @fawfulfan what's been debunked is Hillary's electability. it was fragile &amp; it broke.
Doubting_Tom|vacuumslayer|-0.2714|0.137|0.769|0.093|"@vacuumslayer ""I'm sure *this* tweet about how terrible Hillary and the DNC are will take down Trump once and for all!"""
johnmarkez24|supporthillary|0.508|0.0|0.798|0.202|Show our support for our next president! Hillary for 2016! Click this: https://t.co/UxwV7lmoAL https://t.co/EP1oU7OQAQ
LizardG|qstafford50|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
LizardG|palmerreport|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
Izabelly_paulaa|GirlyofRauhl|-0.5449|0.163|0.837|0.0|RT @GirlyofRauhl: Verdadeiro motivo pela Hillary ter apagado aqueles e-mails! Eram nudes do Justin Bieber! BELIEBERS NO COMANDO #ARIASJUSTI
shitshowdotinfo|katherinejnowak|0.0772|0.104|0.779|0.117|"RT @katherinejnowak: neera has yet to respond with specific errors the dems + hillary's team made; help her out, fam https://t.co/oVuhu75yDS"
shitshowdotinfo|twitter|0.0772|0.104|0.779|0.117|"RT @katherinejnowak: neera has yet to respond with specific errors the dems + hillary's team made; help her out, fam https://t.co/oVuhu75yDS"
grownfairytale|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
farmgurl3|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
Hillary_nataly|_Concubinato|-0.296|0.104|0.896|0.0|"RT @_Concubinato: Alguien ya escucho ""ya no mas"" version acustico de @MicroTDH ? que clases de rap, sos un fenomeno pai"
sbprice|Ian56789|-0.4588|0.13|0.87|0.0|RT @Ian56789: Remember when Russian Hackers forced Hillary to wipe her server after being served with a Congressional Sub Poena to preserve
RaytronixSales|Bryan700|-0.6597|0.265|0.735|0.0|RT @Bryan700: Democrats Attack Donald Trump's Legitimacy After The Baseless Reports Hillary Lost Due to Russian Hackers.
RayneNGrace|dcexaminer|-0.5859|0.232|0.669|0.099|"@dcexaminer Just stop.  Not true.  Hillary is not President because of Hillary, her corruption, the evil in the DNC, the egos.  #FakeNews"
KostJason|JustinRaimondo|-0.8724|0.365|0.635|0.0|"RT @JustinRaimondo: Mr. President, you defeated the media just as you defeated Hillary &amp; they'll never forgive you. Not to worry - your vic"
SusanSt08942260|CronkiteSays|-0.3818|0.205|0.697|0.098|RT @CronkiteSays: REAL NEWSWe've completed an extensive analysis into why Hillary lost and have determined Hillary caused Hillary to lose
constantino_sam|pinterest|-0.8056|0.377|0.623|0.0|DOES THIS ASS MAKE MY TRUCK - ANTI HILLARY PRO TRUMP POLITICAL BUMPER STICKER https://t.co/CZwvohqldH
Mistysmom1|Atrustynote|0.0|0.0|1.0|0.0|RT @Atrustynote: @ANOMALY1 one more time --Hillary Is going back to Arkansas https://t.co/qMNMmtblKG
Mistysmom1|twitter|0.0|0.0|1.0|0.0|RT @Atrustynote: @ANOMALY1 one more time --Hillary Is going back to Arkansas https://t.co/qMNMmtblKG
jopoleski|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
jopoleski|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
KingTurd63|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
aplemkseriously|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
aplemkseriously|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
textifyer59|geordielester|0.4215|0.0|0.872|0.128|"RT @geordielester: russia shouldn't choose the president of the united states. americans should choose, and america chose hillary. this mes"
jjburdett|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
reblor|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
reblor|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
Tymeeks98|tech2eets|-0.3089|0.22|0.78|0.0|@tech2eets @Mitch_John573 Didn't Mexico help Hillary in the election? 
MrJamesonNeat|ArianeBellamar|0.0|0.0|1.0|0.0|RT @ArianeBellamar:  b4 Partisan! Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/CMOS
MrJamesonNeat|t|0.0|0.0|1.0|0.0|RT @ArianeBellamar:  b4 Partisan! Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/CMOS
sandybelyeu|albamonica|0.6124|0.0|0.8|0.2|"RT @albamonica: After the Reid event, Hillary Clinton greeted several Kaine staffers and young supporters, some of whom can be heard sobbin"
fernanda_24680|GirlyofRauhl|-0.5449|0.163|0.837|0.0|RT @GirlyofRauhl: Verdadeiro motivo pela Hillary ter apagado aqueles e-mails! Eram nudes do Justin Bieber! BELIEBERS NO COMANDO #ARIASJUSTI
BTW_LOL|latimes|-0.6971|0.346|0.453|0.201|@latimes NO TIME TO LAUGH. THIS IS SERIOUS. ISIS WILL KILL US ALL. #OBAMA IN HAWAII. #HILLARY LIED TO #FBI... NOT FUNNY AT ALL
SLYBUTCH01|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Sheilas11|mikeoconnor123|-0.7906|0.32|0.68|0.0|"RT @mikeoconnor123: Press said  bi-partisan outrage if Trump challenged election, Then Hillary did just that.  Silence. Story on outrage is"
michele5411|DustinGiebel|-0.4019|0.172|0.828|0.0|RT @DustinGiebel: Hillary hacked the DNC because Trump was hogging all the attention.  #BoltonFalseFlagExcuses
eve1753cm|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
Groughy|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
mimimayesTN|ed_hooley|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
mimimayesTN|truthfeed|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
Britainboy|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
GunnarBj|kpoulsen|-0.7367|0.275|0.725|0.0|"RT @kpoulsen: Icymi, the ""not sure"" part is that Russia's goal may have been to defeat Hillary, not support her opponent https://t.co/2ubio"
GunnarBj|t|-0.7367|0.275|0.725|0.0|"RT @kpoulsen: Icymi, the ""not sure"" part is that Russia's goal may have been to defeat Hillary, not support her opponent https://t.co/2ubio"
Mistysmom1|Atrustynote|0.0|0.0|1.0|0.0|RT @Atrustynote: @ANOMALY1 Hillary's Back Story Is Ghosts Smashed Her Phones &amp; Emails The night Tooth Ferry Visited her home https://t.co/1
Mistysmom1|twitter|0.0|0.0|1.0|0.0|RT @Atrustynote: @ANOMALY1 Hillary's Back Story Is Ghosts Smashed Her Phones &amp; Emails The night Tooth Ferry Visited her home https://t.co/1
breadlightning|katherinejnowak|-0.5267|0.175|0.825|0.0|53. keeping independents out of the primaries made them feel distrusted by Hillary's campaign @katherinejnowak @teeg_dougland @neeratanden
AndreFrato|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
AndreFrato|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
mariemc11308417|LibertyLivesHer|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
mariemc11308417|vivaliberty|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
JayS2629|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
rjber15|WeAreChangeNYC|-0.6124|0.244|0.669|0.087|RT @WeAreChangeNYC: Hillary Clinton Calls For Congress To Go After Fake News Despite Creating Fake News Herself In The Past:https://t.co/
rjber15|t|-0.6124|0.244|0.669|0.087|RT @WeAreChangeNYC: Hillary Clinton Calls For Congress To Go After Fake News Despite Creating Fake News Herself In The Past:https://t.co/
NathanCarreon10|gerfingerpoken|0.0772|0.149|0.683|0.168|RT @gerfingerpoken: Did IRS Leak Trump Returns 2 Help Hillary? https://t.co/EWkqWLPAQNAmerican Thinker https://t.co/L7h6rlr1le https://t.
NathanCarreon10|t|0.0772|0.149|0.683|0.168|RT @gerfingerpoken: Did IRS Leak Trump Returns 2 Help Hillary? https://t.co/EWkqWLPAQNAmerican Thinker https://t.co/L7h6rlr1le https://t.
Catdog2many|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
nobleba|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
AaronHill_|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
serendipity5460|carlbernstein|-0.0477|0.069|0.931|0.0|"@carlbernstein @JoyAnnReid not a single coherent defense of Trump that doesn't start w/ ""but Hillary"" or ""but Obama"" "
CoffeyLiqueur|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
CoffeyLiqueur||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
MisterAK47|brittfpark|-0.4767|0.341|0.659|0.0|RT @brittfpark: Hillary's fake news. #MAGA https://t.co/vbCRiw77D8
MisterAK47|twitter|-0.4767|0.341|0.659|0.0|RT @brittfpark: Hillary's fake news. #MAGA https://t.co/vbCRiw77D8
emccoy_writer|runwithskizzers|0.1603|0.0|0.925|0.075|"RT @runwithskizzers: 500k hearings on Benghazi to confirm that Hillary wasn't at fault, but you won't lift a finger about RUSSIA infiltrati"
SURFER13HB|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
jwire|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
AlirahChristi|KatieWagnerFox|0.3818|0.134|0.634|0.231|"RT @KatieWagnerFox: Seth Rich narc'd DNC emails because of cheating in Primary to promote Hillary. #SethRich, ultimate Bernie Bro, RIP. #"
unixwhisperer|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/T2RfG3mDes via @Change
unixwhisperer|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/T2RfG3mDes via @Change
sliman12|StephensWSJ|0.5719|0.0|0.783|0.217|@StephensWSJ Trump will be much better for Israel than Hillary ever would have been. Bibi agrees 60 minutes tonight.
67purple|ThePatriot143|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
67purple|truthfeed|-0.5319|0.177|0.823|0.0|RT @ThePatriot143: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
MaryhamptonLou|KellyannePolls|0.0|0.0|1.0|0.0|"@KellyannePolls @Newsweek If so, they had rather deal with a man of esteem than dilly dally with crooked Hillary."
catlover1943|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
mikew6161|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
mikew6161||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
MsDemeanor0125|ed_hooley|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
MsDemeanor0125|truthfeed|0.3818|0.0|0.86|0.14|RT @ed_hooley: FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwit
chris63414391|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
mikeman_larson|Snapchat|0.4404|0.0|0.884|0.116|"I feel that if @Snapchat took away the dog filter, there would be more white girls rioting all over the country than Hillary supporters"
nana5greatgrand|ed_hooley|0.0|0.0|1.0|0.0|RT @ed_hooley: DECLINE OF THE DEMOCRATS. JFK SENT MEN TO THE MOON... OBAMA SENT MEN TO THE LADIES ROOM #obama #Hillary #ImWithHer https://t
nana5greatgrand||0.0|0.0|1.0|0.0|RT @ed_hooley: DECLINE OF THE DEMOCRATS. JFK SENT MEN TO THE MOON... OBAMA SENT MEN TO THE LADIES ROOM #obama #Hillary #ImWithHer https://t
marfoglio777|pdachil|0.0|0.0|1.0|0.0|@pdachil @HillaryClinton And Hillary continues to hoard the cash after all the calls for her to return it during election.
JeremyHimli|shoahnuffin1|0.765|0.084|0.617|0.299|@shoahnuffin1 Grow up. You're a big boy. You know better. Hillary is Trump's friend. Always has been. He lied to you a lot. Wise up.
ggbootsrock|charliekirk11|0.0|0.0|1.0|0.0|"RT @charliekirk11: Russia potentially being involved is a big deal, but where was the media when Hillary funded her entire staff with forei"
DesiaAllyJoseph|RepStevenSmith|0.0772|0.0|0.939|0.061|RT @RepStevenSmith: Want to hear about what Hillary did in Libya from a real journalist? @wikileaks Julian Assange explains it in 2 minutes
Dimipace|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
peytonnbrianna|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
PrettyBeaches|ApocalypticaNow|-0.0346|0.077|0.852|0.071|"RT @ApocalypticaNow: I'll never forget how @MSNBC, @CNN &amp; @FoxNews aired an empty podium at a Trump rally instead of a Clinton speech https"
jan5261|peddoc63|-0.5574|0.141|0.859|0.0|RT @peddoc63: Did Russians have anything 2do with DNC &amp; Hillary cheating Bernie out of nomination. Or with media providing Hillary with deb
flajeffreyt|peterdaou|-0.25|0.152|0.738|0.111|"RT @peterdaou: If you're convinced that Hillary is corrupt, flawed, unlikable, dishonest, that was EXACTLY the goal of Russian tampering. C"
TraciGrrl|kylegriffin1|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
TraciGrrl|theatlantic|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
cmgarner_garner|thehill|0.0|0.0|1.0|0.0|"@thehill And Hillary is Mother Teresa, right?"
Benwest2016|LucyAppa|0.0|0.0|1.0|0.0|@LucyAppa @trumpencexual @Salon29Main @CrozieX112 @TerrynRob they always deflect to Hillary.
angelnphx|kurteichenwald|-0.2382|0.22|0.67|0.11|"RT @kurteichenwald: No offense, @chucktodd, but when u say no one was sure Russia behind hack pre-election, shows u need to read more. http"
WendyLynnxoxo|trumpwallnow|0.0|0.0|1.0|0.0|RT @trumpwallnow: I just found what I'm getting Hillary for Christmas. They come in different colors to match her jumpsuits!https://t.co/v
WendyLynnxoxo|abhinavvadrevu|0.0|0.0|1.0|0.0|RT @trumpwallnow: I just found what I'm getting Hillary for Christmas. They come in different colors to match her jumpsuits!https://t.co/v
Debbiemom|Change|0.0|0.0|1.0|0.0|Federal Court: Federal court install Hillary Clinton as POTUS due to Russian Interference in our elec... https://t.co/4c30BCRAsL via @Change
Debbiemom|change|0.0|0.0|1.0|0.0|Federal Court: Federal court install Hillary Clinton as POTUS due to Russian Interference in our elec... https://t.co/4c30BCRAsL via @Change
JEL248|dr2deadline|0.0|0.0|1.0|0.0|@dr2deadline Er det mest relevante ikke at de emails afslrede en korrupt Hillary Clinton? Hvorfor snakkede i ikke om dt? #DKmedier
RamBoPirate|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
7tips1|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
cb55uic|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
hexogennotsugar|thepeoplesview|0.0|0.0|1.0|0.0|RT @thepeoplesview: There are two white men Putin helped in 2016. Both of them ran against Hillary Clinton.
james_towner|FrankLuntz|-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
james_towner||-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
JeremyR1992|Slate|-0.521|0.241|0.669|0.091|"@Slate For some idiotic and strange reason, people won't be alarmed until it somehow lands in Hillary's inbox"
kylorenwashere|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
cfn_ms|lukeoneil47|-0.6597|0.293|0.707|0.0|RT @lukeoneil47: The Democrats hacked the election and emails ...but to make Hillary lose https://t.co/QstENq3dbl
cfn_ms|twitter|-0.6597|0.293|0.707|0.0|RT @lukeoneil47: The Democrats hacked the election and emails ...but to make Hillary lose https://t.co/QstENq3dbl
DoughnutJane|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
JehanneMc|twitter|0.5423|0.0|0.8|0.2|"Yes, my family decided to have Hillary on the top of our Christmas tree this year. #angel #bae #imstillwithher https://t.co/1mA2h546OD"
LAMOONLYNN|bfraser747|-0.6901|0.222|0.778|0.0|"RT @bfraser747:  ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."" ~ @GovMikeHu"
carolinelv|pete03217|-0.8519|0.283|0.717|0.0|RT @pete03217: @lidiya_selwood @suzost @washingtonpost We see it but Dems choose not to see it. They are blind to all the horrible things H
unspokenbond|KatieWagnerFox|0.3818|0.134|0.634|0.231|"RT @KatieWagnerFox: Seth Rich narc'd DNC emails because of cheating in Primary to promote Hillary. #SethRich, ultimate Bernie Bro, RIP. #"
Catdog2many|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
AllNewsDaily|mediaite|0.0|0.0|1.0|0.0|#Breaking #HIllaryNews Former U.S. Ambassador to Russia: Vladimir Putin Wanted 'Revenge' on Hillary Clinton - M... https://t.co/nl5QVak8mD
crkienast|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
andrewfriedman0|DrJillStein|0.0258|0.2|0.596|0.204|"@DrJillStein Yep, no difference in Trump and Hillary. Except on Choice. Immigration. Unions. Supreme Court. Minimum Wage. Etc. Fuck You Jill"
Black_Feather55|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
clintonistaa|HillaryTheBOSS|0.0|0.0|1.0|0.0|RT @HillaryTheBOSS: Hillary del Rodman  https://t.co/O5aanBZoQd
clintonistaa|twitter|0.0|0.0|1.0|0.0|RT @HillaryTheBOSS: Hillary del Rodman  https://t.co/O5aanBZoQd
alpaca500|GarbageTime01|0.0|0.0|1.0|0.0|"RT @GarbageTime01: @PussyGrabber45 @KellyannePolls @nypost Hillary's campaign was funded by Saudi Arabia. And thats proven, unlike the Russ"
LiftedTitan|bessbell|-0.7089|0.228|0.772|0.0|"@bessbell @realDonaldTrump By the way, Hillary was proven guilty of having a private very insecure server. You know why they let her off?"
Zina_Solomon|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 https://t.co/6GnySGv9eR via @Change
Zina_Solomon|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 https://t.co/6GnySGv9eR via @Change
johnsenrm|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
genyorke|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
badger3030|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
1isten_up|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
LizalcornLiz|ed_hooley|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
LizalcornLiz|truthfeed|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
ggbootsrock|ed_hooley|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
ggbootsrock|truthfeed|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
jsirwin67|blackagendareport|-0.743|0.441|0.559|0.0|"Libya: Hillarys War, the Empires Mistake | Black Agenda Report https://t.co/7p7FrECrI5"
gerfingerpoken|IBDeditorials|0.431|0.0|0.82|0.18|(IBD) Hillary Rodham Nixon - Even He Didn't Destroy The Tapes  - https://t.co/OnpEFahSgW - @IBDeditorials - https://t.co/RCL5K0tY1i 11
gerfingerpoken|investors|0.431|0.0|0.82|0.18|(IBD) Hillary Rodham Nixon - Even He Didn't Destroy The Tapes  - https://t.co/OnpEFahSgW - @IBDeditorials - https://t.co/RCL5K0tY1i 11
SheilaDecker19|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
brenny_|RNRMississippi|-0.2263|0.215|0.642|0.143|"RT @RNRMississippi: Russians are Amazing: Set up a private server, rigged the primary, used BleachBit to violate a court order, then made"
JSavoly|addictinginfo|-0.7378|0.342|0.658|0.0|Silvers Election Autopsy And Reason For Hillarys Loss Will INFURIATE Everyone #StollenElection #ComradeTrump  https://t.co/vpyHU4Ts6n
k_brucks|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
silver_selkie|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
silver_selkie|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
leameadow|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
78izzie|ed_hooley|-0.7269|0.337|0.663|0.0|RT @ed_hooley: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/RKOyB0S2vR
78izzie|nytimes|-0.7269|0.337|0.663|0.0|RT @ed_hooley: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/RKOyB0S2vR
MiaEvan30311368|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
Gan1Nancy|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
MissSweets2|ed_hooley|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
MissSweets2|truthfeed|0.0|0.0|1.0|0.0|"RT @ed_hooley: British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
phred47|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
JoyPuder|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
Bugsben20|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
OatesTuzzio|HuffingtonPost|-0.7506|0.252|0.748|0.0|@HuffingtonPost sadly many bitched that Hillary had the nerve 2 wear pants. Sexist. Even some women. But new hashtag for cabinet #ToxicWaste
divadarya|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
RalphHornsby|americanlookout|0.0|0.0|1.0|0.0|Morning Joes Mika: The Hillary Clinton Campaign Wanted Me Pulled Off The Air (VIDEO)  American Lookout https://t.co/ODpj9gwtNR
gpnavonod|GodandtheBear|-0.8225|0.388|0.612|0.0|"RT @GodandtheBear: Hillary is the worst of bad people, a wolf in sheep's clothing. https://t.co/wy3ux6sLx9"
gpnavonod|twitter|-0.8225|0.388|0.612|0.0|"RT @GodandtheBear: Hillary is the worst of bad people, a wolf in sheep's clothing. https://t.co/wy3ux6sLx9"
mildredshackle1|Humans_vs_Trump|0.34|0.099|0.719|0.182|RT @Humans_vs_Trump: Hillary Clinton hates the spotlight &amp; likes doing the work. Imagine what it must be like for her to read headline. htt
egopanthers|NateSilver538|-0.3182|0.103|0.897|0.0|"@NateSilver538 Hillary Clinton had the biggest impact on the election, she blew $1 1/4 Bllion and still lost b/c sh https://t.co/BPYxBqt0FJ"
egopanthers|twitter|-0.3182|0.103|0.897|0.0|"@NateSilver538 Hillary Clinton had the biggest impact on the election, she blew $1 1/4 Bllion and still lost b/c sh https://t.co/BPYxBqt0FJ"
ThatGuyMelts|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
ThatGuyMelts|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
MyCrashIs|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
syqau|syqau|-0.6351|0.224|0.776|0.0|"RT @syqau: During recount, in 100 precincts in Milwaukee, WI,  Hillary Clinton lost 17,000 votes!! (Trump lost only 1,700) https://t.co/VS"
syqau|t|-0.6351|0.224|0.776|0.0|"RT @syqau: During recount, in 100 precincts in Milwaukee, WI,  Hillary Clinton lost 17,000 votes!! (Trump lost only 1,700) https://t.co/VS"
whitemomgoals|LifeWinnersOnly|-0.6124|0.278|0.722|0.0|RT @LifeWinnersOnly: Hillary Campaign Ignored Staffer Who Predicted She'd Lose | The Daily Caller https://t.co/VEWulSEspS #breaking
whitemomgoals|dailycaller|-0.6124|0.278|0.722|0.0|RT @LifeWinnersOnly: Hillary Campaign Ignored Staffer Who Predicted She'd Lose | The Daily Caller https://t.co/VEWulSEspS #breaking
miller_jeneal|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
bloodinbritish3|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
marieann66|rodimusprime|0.4019|0.0|0.856|0.144|"@rodimusprime @EmilyWhiteUSA1 Yes, the Independent Sanders that along with GOP helped elect Trump with his Hillary trashing."
frodofied|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
roqchrisy|kimconde752|0.0|0.0|1.0|0.0|RT @kimconde752: #meetthepress @chucktodd @AdamSchiffCA explain how Hillary Clinton stood up to the Russians? Was before or after she sold
jmingerson725|Sherrishaw14|0.0|0.0|1.0|0.0|RT @Sherrishaw14: @whirrll @FredPecora @GOP @PatriotsOfMars @freep Hillary is the only one who can finish this https://t.co/uoRiqedjhA
jmingerson725|twitter|0.0|0.0|1.0|0.0|RT @Sherrishaw14: @whirrll @FredPecora @GOP @PatriotsOfMars @freep Hillary is the only one who can finish this https://t.co/uoRiqedjhA
rowilkins|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
ldiproperzio|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
winkiechance|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
MyPupVoted|JustNWashington|0.0|0.0|1.0|0.0|RT @JustNWashington: Hillary's response to a reporter asking her if she'd ever lied... https://t.co/dmVw3IvoYq
MyPupVoted|twitter|0.0|0.0|1.0|0.0|RT @JustNWashington: Hillary's response to a reporter asking her if she'd ever lied... https://t.co/dmVw3IvoYq
SamWiseMD|Dan_Roehm|0.0|0.0|1.0|0.0|"RT @Dan_Roehm: the map of the leftist Hillary majority vs the ""minority"" of all American votes really tells a story. 98% of the US land mas"
ChaosApathy|SLindauer2011|-0.2808|0.178|0.697|0.125|RT @SLindauer2011: QUEEN OF FAKE NEWS: 8 Times Hillary Fabricated Stories to Help Her Image https://t.co/fKGb8D3RfS via @regisgiles
ChaosApathy|girlsjustwannahaveguns|-0.2808|0.178|0.697|0.125|RT @SLindauer2011: QUEEN OF FAKE NEWS: 8 Times Hillary Fabricated Stories to Help Her Image https://t.co/fKGb8D3RfS via @regisgiles
MstrWaterbender|HumanistReport|-0.25|0.156|0.769|0.075|"RT @HumanistReport: Hillary Clinton split the party, moved liberals to the right, and normalized war mongering, but still claims to be the"
JBVenn|dandrezner|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
JBVenn|t|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
paulbenedict7|paulbenedict7|-0.7906|0.333|0.667|0.0|RT @paulbenedict7: #Obamastan's FBI: no need to prosecute Hillary's uranium deal; Obamastan's CIA: Putin is a #Trump lobbyist. Worse than #
Quicksilver2723|theGSpledge|0.0|0.0|1.0|0.0|"RT @theGSpledge: If there's 1 thing Hillary's disappearance in the face of Trump shows is that she never was a leader, just a self-entitled"
Tuigen|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
meatball_writes|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
VCooper51|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
AliBakirdan|twitter|0.4588|0.0|0.85|0.15|I am glad to see that Hillary Clinton has a hashtag trending about her heavy use of medications. #married2med https://t.co/L2MN3E1Sce
Col_Connaughton|youtube|-0.2003|0.121|0.879|0.0|Fox News Exposes George Soros &amp; Hillary Clinton Relationship! https://t.co/NCVoB6NemR #hillary #clinton #soros #BLM
janiceponchak|cramer_here|0.0|0.0|1.0|0.0|RT @cramer_here: #TRUMP WON!#HILLARY LOST!#my4wordfails
Buiock|BreezeCyclone|0.3802|0.0|0.868|0.132|@BreezeCyclone @TayTay78730804 By kicking Hillary out world  dodged a huge bullet .On same Level as Sharia or the Nazis!
SaltSashi|kylegriffin1|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
SaltSashi|theatlantic|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
TheOneLadyEagle|ReversingASD|0.0|0.0|1.0|0.0|RT @ReversingASD: Fox News LiveHILLARY BELONGS IN JAIL! TREY GOWDY VS HILLARY CLINTON US News Today https://t.co/tuqjfyKmNF via @youtube
TheOneLadyEagle|youtube|0.0|0.0|1.0|0.0|RT @ReversingASD: Fox News LiveHILLARY BELONGS IN JAIL! TREY GOWDY VS HILLARY CLINTON US News Today https://t.co/tuqjfyKmNF via @youtube
kingvideo123|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
Psychotic_Beast|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 https://t.co/JyKhUGriA9 via @Change
Psychotic_Beast|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 https://t.co/JyKhUGriA9 via @Change
nauthizjane|thehill|-0.3818|0.115|0.885|0.0|Bolton has a point. How  many times have Obama and Hillary lied to us? How many times has Obama used the... https://t.co/TX3tCKC8KX
DCoryReynolds|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
syqau|syqau|-0.128|0.13|0.87|0.0|RT @syqau: Alcoholism has contributed to Hillary Clinton's lowered IQ... https://t.co/dxd7hHyqOl
syqau|twitter|-0.128|0.13|0.87|0.0|RT @syqau: Alcoholism has contributed to Hillary Clinton's lowered IQ... https://t.co/dxd7hHyqOl
SscottSsmith84|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
DennisKulpa|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
DennisKulpa||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
Trues55|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
ModernDayZorro|Wikileaks|-0.3818|0.178|0.822|0.0|Fox News FBI @Wikileaks just took a dump on hillary clinton: https://t.co/SLqPGbcxeh via @YouTube
ModernDayZorro|youtube|-0.3818|0.178|0.822|0.0|Fox News FBI @Wikileaks just took a dump on hillary clinton: https://t.co/SLqPGbcxeh via @YouTube
caroljdavy|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @PosyBass1 @SocialCivility it means that in Racine, as votes were counted, Hillary Clinton's large percentage declined +"
ModernDayZorro|YouTube|-0.4767|0.181|0.819|0.0|"HILLARY CLINTON COST HILLARY CLINTON THE ELECTION, Not Fake News Joe Scarborough: https://t.co/V304n1KiSB via @YouTube"
ModernDayZorro|youtube|-0.4767|0.181|0.819|0.0|"HILLARY CLINTON COST HILLARY CLINTON THE ELECTION, Not Fake News Joe Scarborough: https://t.co/V304n1KiSB via @YouTube"
HartmanSeth14|ConservativeFB|-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
HartmanSeth14||-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
ModernDayZorro|YouTube|-0.1531|0.191|0.648|0.161|FOX NEWS FBI READY TO INDICT HILLARY EVIDENCE 'WORSE THAN ANYONE THINKS: https://t.co/8CNGPeeJ3S via @YouTube
ModernDayZorro|youtube|-0.1531|0.191|0.648|0.161|FOX NEWS FBI READY TO INDICT HILLARY EVIDENCE 'WORSE THAN ANYONE THINKS: https://t.co/8CNGPeeJ3S via @YouTube
darlingrue|peterdaou|-0.0173|0.128|0.746|0.126|"RT @peterdaou: TRUTH: Hillary's ""unlikability"" WAS the Russian strategy. Make her toxic with fake news, trolling, hacking. 66 million didn"
ancerrone|CarmineZozzora|0.85|0.0|0.634|0.366|RT @CarmineZozzora: Russian hacking narrative mysteriously absent when Hillary was sure to win - but magically surfaces after Trump's win?
Byrlyne|bfraser747|-0.6901|0.222|0.778|0.0|"RT @bfraser747:  ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."" ~ @GovMikeHu"
AllNewsDaily|mediaite|0.0|0.0|1.0|0.0|#ShesWithUs | Former U.S. Ambassador to Russia: Vladimir Putin Wanted 'Revenge' on Hillary Clinton - Mediaite https://t.co/lxkAp3Ndao
KenEhrhart|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
KenEhrhart|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
Ethan115x|RealDonaldTurn|0.5719|0.0|0.448|0.552|@RealDonaldTurn @Chaosxsilencer Hillary won
COS_PalmBayFL|ambitjournal|-0.128|0.254|0.563|0.183|RT @ambitjournal: Hillary loved fake news  until she lost | Guest Column | World | News | Toronto https://t.co/z3T8xDO2YT
COS_PalmBayFL|torontosun|-0.128|0.254|0.563|0.183|RT @ambitjournal: Hillary loved fake news  until she lost | Guest Column | World | News | Toronto https://t.co/z3T8xDO2YT
Avg_Voter|BrittPettibone|-0.8316|0.468|0.532|0.0|RT @BrittPettibone: Kellyanne Conway is battling a barrage of death threats from Hillary Supporters.#FridayFeelinghttps://t.co/0kLbme7ouQ
Mcatlady54|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
HollyCarolEarls|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
HollyCarolEarls|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
courthulsart|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
ZarkoElDiablo|DarinDorsey4|-0.4512|0.176|0.745|0.079|RT @DarinDorsey4: @mitchellvii @ZarkoElDiablo @HillaryClinton I rarely disagree will @mitchellvii but the problem with Hillary was she was
linos2015|HispanicsTrump|0.7579|0.0|0.764|0.236|RT @HispanicsTrump: Sometimes it's nice to just sit back and be thankful that Hillary Clinton won't be our next president. Everything is lo
pkhinkle|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
ukexpat19|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
ukexpat19|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
TiffanieAnn16|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
DavidLance3|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Millenniumistic|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/1zCwaCuFYY via @Change
Millenniumistic|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/1zCwaCuFYY via @Change
monkeynaut1966|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
_StarlightLive_|octaviahenke|-0.5719|0.236|0.647|0.117|"RT @octaviahenke: @FoxNews Obama needs to pack his things and get ready to get out, your flunky Hillary lost. Its over. No matter what you"
ThreatcoreNews|smerconish|-0.4019|0.252|0.748|0.0|.@smerconish I guess the Russians hacked Hillary's crowds too? #investigate
mrchristopher03|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
mrchristopher03|t|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
geoff_deweaver|DRUDGE_REPORT|-0.5574|0.217|0.783|0.0|RT @DRUDGE_REPORT: Madonna and Hillary: 'Witch' and 'Nasty Woman' as Sisters in Arms... https://t.co/htlaxNPgSe
geoff_deweaver|nytimes|-0.5574|0.217|0.783|0.0|RT @DRUDGE_REPORT: Madonna and Hillary: 'Witch' and 'Nasty Woman' as Sisters in Arms... https://t.co/htlaxNPgSe
wheelchairant|imfsea_aruna|-0.2263|0.164|0.711|0.124|@imfsea_aruna @DrJillStein @Cosmopolitan Most likely did with Hillary's popular vote and his anger over recounting which is constitutional.
victor81054|MikaelaSkyeSays|-0.296|0.121|0.879|0.0|RT @MikaelaSkyeSays: @jilevin - And the media refused to cover this.  But Hillary's deplorable comment got 24/7 coverage.
ed_hooley|truthfeed|0.3818|0.0|0.843|0.157|FLASHBACK VIDEO : Obama Busted on HOT MIC Making Secret Promises Russia https://t.co/thZymgbdUS#maga #obama #hillary #imwithher
1sfleming302|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: People weren't concerned about Russia when Hillary was selling them US uranium.#MAGA
SoapView|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
AugustusFaber|RNRMississippi|-0.2263|0.215|0.642|0.143|"RT @RNRMississippi: Russians are Amazing: Set up a private server, rigged the primary, used BleachBit to violate a court order, then made"
FergKei|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
FergKei|t|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
heatherduffer|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
pjmcgovern4|Im_ConnorKelley|0.5719|0.0|0.73|0.27|RT @Im_ConnorKelley: @realDonaldTrump @NBCNightlyNews @CNN Hillary won by 2.83 million votes
tangytangier|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
Gan1Nancy|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
Gan1Nancy|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
bourgeoisalien|realDonaldTrump|0.7221|0.127|0.559|0.315|@realDonaldTrump  @CNN congrats on requesting clearance for a conspiracy nut who claims Hillary operates a Satanic child-sex ring! SO SMART!
FisherBurton|BillyVonElds|-0.5994|0.243|0.681|0.077|"@BillyVonElds No, anyone who sees that is fine with Hillary's pro-fracking, pro-pipeline, pro-wall St. warmongering and really blew it."
Freedom1776__|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
LoveOireachtas|halsteadg048|0.0|0.0|1.0|0.0|RT @halsteadg048: Hillary Clinton Takeover of the USA https://t.co/WyvI6OVBrT PROOF By Dr Pieczenik Counter-Coup Who Worked w/ Julian To St
LoveOireachtas|youtube|0.0|0.0|1.0|0.0|RT @halsteadg048: Hillary Clinton Takeover of the USA https://t.co/WyvI6OVBrT PROOF By Dr Pieczenik Counter-Coup Who Worked w/ Julian To St
StormSpinning|DisabilityPower|-0.3716|0.124|0.876|0.0|"RT @DisabilityPower: @womensmarch I march because Hillary took on Russia, FBI, white supremecy, Ableism, Racism &amp; Sexism; but never gave u"
lkmcland|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
lkmcland||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
MissEMT37|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
123andgo|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
deorhtayxkvwmp1|sexdatehere2|0.0|0.0|1.0|0.0|teen hillary scottcurry https://t.co/ANhGjtKcKs
1isten_up|guntrust|0.0|0.0|1.0|0.0|RT @guntrust: Wikileaks: Dana Loesch - Hillary's Middle Eastern Firearms Deals Sent Cash to Clinton https://t.co/QVYT2lZhGR #tcot #ccot #2A
1isten_up|lawnews|0.0|0.0|1.0|0.0|RT @guntrust: Wikileaks: Dana Loesch - Hillary's Middle Eastern Firearms Deals Sent Cash to Clinton https://t.co/QVYT2lZhGR #tcot #ccot #2A
MarkShawnda|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
FlippinDBird|BrotherVet|0.6037|0.0|0.753|0.247|RT @BrotherVet: @RoyalTXGirl @sharon4marie @FlippinDBird @940heidiWONDER IF HILLARYS DONOR CARE https://t.co/BEshBi0nE7 via @dailycaller
FlippinDBird|linkis|0.6037|0.0|0.753|0.247|RT @BrotherVet: @RoyalTXGirl @sharon4marie @FlippinDBird @940heidiWONDER IF HILLARYS DONOR CARE https://t.co/BEshBi0nE7 via @dailycaller
bpman1973|Cernovich|0.296|0.083|0.795|0.123|"RT @Cernovich: If Hillary had won we'd have talked about ""rigged elections"" for a day or two and then moved on. What we are seeing today is"
palestininianpr|MaxBlumenthal|0.0|0.0|1.0|0.0|RT @MaxBlumenthal: .@AliAbunimah @JoyAnnReid What we've learned here is that Putin took out Hillary but Hillary did not take out Qaddafi. h
ReginaPeele|albamonica|0.6124|0.0|0.8|0.2|"RT @albamonica: After the Reid event, Hillary Clinton greeted several Kaine staffers and young supporters, some of whom can be heard sobbin"
NotouriosJew|ifunny|0.0|0.0|1.0|0.0|#hillary #hillaryclinton #election #trumpadministration #trump https://t.co/l7QDtK5lnx https://t.co/XbTnvUf7mT
bigdieseldan04|SamanthaClarkH|-0.4824|0.164|0.836|0.0|"RT @SamanthaClarkH: FBI ASST. DIRECTOR COMES OUT, Says HILLARY SHOULD BE SHOT BY FIRING SQUAD https://t.co/HopZEh35Uo https://t.co/e1TInK"
bigdieseldan04|conservativefighters|-0.4824|0.164|0.836|0.0|"RT @SamanthaClarkH: FBI ASST. DIRECTOR COMES OUT, Says HILLARY SHOULD BE SHOT BY FIRING SQUAD https://t.co/HopZEh35Uo https://t.co/e1TInK"
YaPasdePRESSE|yapasdpresse|0.0|0.0|1.0|0.0|#cybercrime Russie ou autres: les Dmocrates responsables des vols de donnes (les choix d'Hillary Clinton) https://t.co/VJu3QKhK32
carolinelv|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
carolinelv|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
Dovemom77|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
sarahsophief|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
joyhaler|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Lancelot_R_King|PARISDENNARD|0.0|0.0|1.0|0.0|RT @PARISDENNARD: JFK had his brother as AG and Hillary Clinton took on policy with an office in the West Wing so it's not uncommon to have
ShaftonP|gerfingerpoken|0.0772|0.149|0.683|0.168|RT @gerfingerpoken: Did IRS Leak Trump Returns 2 Help Hillary? https://t.co/EWkqWLPAQNAmerican Thinker https://t.co/L7h6rlr1le https://t.
ShaftonP|t|0.0772|0.149|0.683|0.168|RT @gerfingerpoken: Did IRS Leak Trump Returns 2 Help Hillary? https://t.co/EWkqWLPAQNAmerican Thinker https://t.co/L7h6rlr1le https://t.
wendellshaw5|S1776frdm|-0.9186|0.519|0.417|0.064|"RT @S1776frdm: Hillary Sucked at everything except Treason Corruption Pay4PlayKindness of Spirit Racism, Hate 4 Average Citizens--https:/"
wendellshaw5||-0.9186|0.519|0.417|0.064|"RT @S1776frdm: Hillary Sucked at everything except Treason Corruption Pay4PlayKindness of Spirit Racism, Hate 4 Average Citizens--https:/"
crkienast|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
bugsy159|Dr_of_Nursing|0.6124|0.0|0.762|0.238|"RT @Dr_of_Nursing: #Treason disqualifies #Trump from being PEOTUS, #ElectoralCollege can easily resolve the issue by choosing #Hillary http"
ThePatriot143|truthfeed|-0.5319|0.197|0.803|0.0|This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House  TruthFeed https://t.co/snLNt7H5W3
2sumextent|CuckStomper|0.1901|0.191|0.629|0.18|"@CuckStomper @RubinReport no, but glad Hillary and her itchy trigger finger is now in the rearview mirror"
TPD1990|DemocratCespool|-0.4939|0.158|0.842|0.0|RT @DemocratCespool: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #clintonfoundation http
kfredrick15|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
TuxiTix4|nyinvesting|0.0|0.0|1.0|0.0|RT @nyinvesting: @America_1st_ @StupidBoomers @GovMikeHuckabee Russians didn't make Hillary go to coal country and say coal workers should
beth_deitchman|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
constantino_sam|pinterest|0.4404|0.0|0.775|0.225|Vote for Monica Lewinsky's Ex-Boyfriend's Wife  Funny Hillary Clinton Anti-Hilla https://t.co/ZAf33aLWGv
honorverity|redwardprice719|-0.228|0.173|0.693|0.134|"RT @redwardprice719: @Khanoisseur @theonlyadult Hillary's said it and it's absolutely true, therefore That Racist is an Illegitimate Presid"
Tturedraider123|FOLLOW_DA_BUCKS|0.4215|0.0|0.843|0.157|RT @FOLLOW_DA_BUCKS: The Hillary Clinton Takeover of the United States  @sharpfang @Goddess300 @RealAlexJones @Deplorarable_Oz Seen thisht
cassidyphoenyx|JustinRaimondo|-0.8724|0.365|0.635|0.0|"RT @JustinRaimondo: Mr. President, you defeated the media just as you defeated Hillary &amp; they'll never forgive you. Not to worry - your vic"
hartsigns|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
IndeCardio|Dan_Roehm|0.0|0.0|1.0|0.0|"RT @Dan_Roehm: the map of the leftist Hillary majority vs the ""minority"" of all American votes really tells a story. 98% of the US land mas"
jacobspm|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
bastiongray|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
rehmanursami|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
linos2015|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
linos2015||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
JackRoss061485|EricKleefeld|0.0|0.0|1.0|0.0|@EricKleefeld An accurate description of what Hillary's position vis-a-vis the Saudis would have been.
LeAnne_Watrous|twitter|0.0|0.0|1.0|0.0|They just can't wrap their brains around the fact that American voters actually wanted Trump over Hillary. https://t.co/EKZIOksMxG
MEUDEUSDOCELL|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
lobaoeletrico|brasil_fotos|0.6124|0.0|0.75|0.25|RT @brasil_fotos: @SV99999 @lobaoeletrico The biggest supporter for ISIS is the main one for Hillary. Funny thing...
bawlaw99|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
bawlaw99|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
starlady24|CapitalismCures|-0.6289|0.293|0.557|0.15|RT @CapitalismCures: Leftists are trying to blame the election results on white supremacy. WRONG. Its because no one trusts Hillary. #Liber
AshPoliceReddy|SpeakerRyan|0.0258|0.11|0.776|0.114|@SpeakerRyan seemed to be eager to speak about Hillary Clinton. Why the reluctance with Donald Trump? Partisan poli https://t.co/iL2n9d459t
AshPoliceReddy|twitter|0.0258|0.11|0.776|0.114|@SpeakerRyan seemed to be eager to speak about Hillary Clinton. Why the reluctance with Donald Trump? Partisan poli https://t.co/iL2n9d459t
AW2B12|jayeljac|-0.5255|0.22|0.78|0.0|@jayeljac @kurteichenwald While they covered Hillary's emails for weeks and months...they ruined Hillary!
THEdavidharris|secureworks|0.0|0.0|1.0|0.0|And SecureWorks added a third independent investigation https://t.co/O13i5ERaO5
agueros_henry|BrittPettibone|0.4404|0.0|0.861|0.139|"RT @BrittPettibone: #ImStillNotOver the fact that, based on zero evidence, Hillary Supporters insist that Russian Hackers interfered in the"
carlettedup|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
miller_jeneal|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: Hillary's secret $2.35M Russian Connection was so crooked, even the #CorruptMedia had to covered it. #UraniumOnehttps://t."
TuxiTix4|willhoerter|0.4755|0.099|0.703|0.197|RT @willhoerter: @America_1st_ @GovMikeHuckabee HILLARY SUCKS EVERYBODY KNOWS THAT BUT THE LITTLE d party still stands for DENIAL.
Coreybez1|WillettKat|-0.5994|0.221|0.692|0.087|RT @WillettKat: Bernies first issue was to destroy Hillary Clinton. He's a traitor to the cause and now just blathers on like a fool about
julainestone|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
julainestone||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
Nessawbu|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
2qris1|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
2qris1|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
FootballKig|TeamTrumpCO|0.0|0.0|1.0|0.0|RT @TeamTrumpCO: #Putin informing #Hillary how he's rigging election!#JillStein=#SCAM#DemocratParty=#Meltdown=#RIP#voterfraud=no #voterI
Phoenixwmn|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: Think bout this: Allied intel servives investigating prez-elect 2 learn if he's Putin stooge in place 2 shatter NATO ht
Skonialo|CindiLewis9|0.1531|0.099|0.776|0.125|"@CindiLewis9 @lives2write4tv You guys need better coping skills. Hillary lost 84% of US counties bc she's an unlikeable, corrupt has-been."
BellaLibelle|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
BellaLibelle|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
antilamegame|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
Zelidasquare|larrywilbur71|-0.4019|0.13|0.87|0.0|"@larrywilbur71 Not machines,they're saying the DNC emails were hacked by Russia and the emails negatively influenced election w/ Hillary"
alllibertynews|tom_tsetung|-0.6023|0.285|0.622|0.093|"RT @tom_tsetung: @Judgenap : Russian didn't hack DNC. The NSA hacked the DNC, bcz they didn't want Hillary, a national security criminal, t"
thefiffer|anylaurie16|0.0|0.0|1.0|0.0|"RT @anylaurie16: President-elect Hillary Clinton gave cabinet positions to 6 major donors, which is unprecedented. https://t.co/MfkBotM6jJ"
thefiffer|twitter|0.0|0.0|1.0|0.0|"RT @anylaurie16: President-elect Hillary Clinton gave cabinet positions to 6 major donors, which is unprecedented. https://t.co/MfkBotM6jJ"
jamesmurphypdx|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
FILLMOE4LIFE|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/s6QHBI9irN via @Change
FILLMOE4LIFE|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/s6QHBI9irN via @Change
rwcox75|anythingbutdem|-0.6808|0.286|0.714|0.0|@anythingbutdem both sides used fake news. But Hillary's team witch was most media ran a lot more
JBax52|DustinGiebel|-0.4019|0.172|0.828|0.0|RT @DustinGiebel: Hillary hacked the DNC because Trump was hogging all the attention.  #BoltonFalseFlagExcuses
bbeaty32|twitter|0.0|0.0|1.0|0.0|"That's nor hillary,  double  https://t.co/NDK0FFhm3w"
jsirwin67|HuffPostPol|-0.5574|0.205|0.795|0.0|"A Vote For Hillary Clinton Is A Vote For Wars Against Russia, China, Others https://t.co/2XAn5aXsK3 via @HuffPostPol"
jsirwin67|huffingtonpost|-0.5574|0.205|0.795|0.0|"A Vote For Hillary Clinton Is A Vote For Wars Against Russia, China, Others https://t.co/2XAn5aXsK3 via @HuffPostPol"
MikeyBong1|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
MWatts08|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
WombatWithWings|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
DavidTravillia1|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
springerpappy|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
ciji2016|peddoc63|0.1531|0.169|0.642|0.189|RT @peddoc63: Hillary left herself vulnerable to hacking &amp; put National Security in jeopardy. Do you care That Obama tried to influence Isr
roqchrisy|NoahBerhe|0.0|0.0|1.0|0.0|RT @NoahBerhe: @RexHuppke Hillary also funded by Saudi government
virleehol|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
anjaligupta90|mitchellvii|0.0|0.0|1.0|0.0|@mitchellvii Dog ate Hillary ballots.
batgirline|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
silverhardt|scottienhughes|-0.8374|0.344|0.656|0.0|@scottienhughes his cabinet choices are the Elitists wasn't that his &amp; all of you liars moaned about with Hillary LIARS
judith_hillary|CrlosElizondo|-0.296|0.239|0.761|0.0|RT @CrlosElizondo: Cuando aplicas sarcasmo y no entienden https://t.co/zj1dpIyg3z
judith_hillary|twitter|-0.296|0.239|0.761|0.0|RT @CrlosElizondo: Cuando aplicas sarcasmo y no entienden https://t.co/zj1dpIyg3z
SscottSsmith84|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
sleepywhiner|twitter|-0.4019|0.351|0.649|0.0|Obama wanted Hillary to lose? https://t.co/fosObs31vw
timtincher|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
ArthurCSchaper|unsavoryagents|0.7506|0.0|0.795|0.205|RT @unsavoryagents: THE DEMOCRATS ARE SO CONCERNED ABOUT RUSSIANS HACKING US BUT DON'T SEEM TO CARE THAT HILLARY HAD A STATE DEPARTMENT SER
NCbgirl|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
JhonRiddik|ebay|0.0|0.0|1.0|0.0|#ChristmasIdeas  Boys Club #1 FIRST APPEARANCE OF PEPE THE FROG Teenage Dinosaur 2006 NM HILLARY https://t.co/Dx3kXPP95S
TravisRuger|kimberlymontse1|0.0|0.0|1.0|0.0|RT @kimberlymontse1: @standupgyrl @TravisRuger as if Hillary's choices would be any different #HelloOligarchy
loriboud|twitter|-0.2023|0.148|0.734|0.119|He is a PATHOLOGICAL LIAR JUST LIKE HILLARY &amp; HES NOT AMERICAN. THEY SAID IMPEACH HIM IN 2011 don't know why they d https://t.co/ldjGYACw4X
notthatCate|dandrezner|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
notthatCate|t|0.6705|0.0|0.776|0.224|"RT @dandrezner: Thank goodness Hillary Clinton, who would have been in the pocket of the donor class, won't be president. https://t.co/8Xx3"
_premiumfan|dashing_reaver|-0.5267|0.195|0.805|0.0|"@dashing_reaver @BillNemacheck ah, Trump is a private citizen, Hillary is a government employee you retard, big difference"
rob_strifeheart|katherinejnowak|0.0772|0.104|0.779|0.117|"RT @katherinejnowak: neera has yet to respond with specific errors the dems + hillary's team made; help her out, fam https://t.co/oVuhu75yDS"
rob_strifeheart|twitter|0.0772|0.104|0.779|0.117|"RT @katherinejnowak: neera has yet to respond with specific errors the dems + hillary's team made; help her out, fam https://t.co/oVuhu75yDS"
MencheyKathleen|c0nvey|0.0|0.0|1.0|0.0|Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted... https://t.co/XRDzA7wBEF by #DailyCaller via @c0nvey
MencheyKathleen|linkis|0.0|0.0|1.0|0.0|Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted... https://t.co/XRDzA7wBEF by #DailyCaller via @c0nvey
travelanita|foxandfriends|0.4019|0.0|0.881|0.119|"@foxandfriends Yes why were Hillary's buddies who she sold US Uranium to, allowing hackers to hack US? If it was Russians"
twolittlestars|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
mariemc11308417|ConservativeFB|-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
mariemc11308417||-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
TuxiTix4|America_1st_|-0.6901|0.222|0.778|0.0|"RT @America_1st_: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candi"
dansheehan|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
dansheehan||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
Cheerful_7|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
reynolds60492|BrowningMachine|-0.3612|0.164|0.746|0.09|@BrowningMachine @Evan_McMullin @realDonaldTrump important to remember mcmuffin was a CIA plant to throw election to Hillary. They failed.
vtgirlinor|npr|0.3612|0.0|0.889|0.111|"U.S. Kids Far Less Likely To Out-Earn Their Parents, As Inequality Grows we can thank Hillary and Trump for this https://t.co/UjCOPjCqUN"
phil4gop|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
dcfodder|fossyboots|0.2944|0.0|0.909|0.091|@fossyboots @Kelebration It was #Hillary who sold 20% of our uranium 2 #Russia and #obama who said he would be more flexible after election
FeistyTrumpette|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
jakesCove_US|trumpwallnow|0.0|0.0|1.0|0.0|RT @trumpwallnow: I just found what I'm getting Hillary for Christmas. They come in different colors to match her jumpsuits!https://t.co/v
jakesCove_US|abhinavvadrevu|0.0|0.0|1.0|0.0|RT @trumpwallnow: I just found what I'm getting Hillary for Christmas. They come in different colors to match her jumpsuits!https://t.co/v
CarlNyberg312|ggreenwald|-0.4588|0.12|0.88|0.0|"I recall GOP/NRA attacking Hillary as too far to the Left on one issue: guns, the one issue where HRC ran to Bernie's Left.@ggreenwald"
salrizzo5|LisaToddSutton|0.7717|0.108|0.518|0.375|@LisaToddSutton @KellyannePolls right she won what's the problem with Hillary lovers to face the truth grow up
skirtyboots|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
Ruthperricone|ConservativeFB|-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
Ruthperricone||-0.4939|0.158|0.842|0.0|RT @ConservativeFB: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #ClintonCash https://t.c
Byrlyne|LVNancy|0.5719|0.0|0.791|0.209|"RT @LVNancy: #RussianHackers IF sore-Loser, Hillary had won, would we be having this conversation?#SundayMorning #TRUMP#AmericaFirst"
Betterw05759703|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: @AchaPatricia You didnt read a lot of what I wrote pre-election, did you? Try these:https://t.co/JSN8Liptfchttps://t."
Betterw05759703|t|0.0|0.0|1.0|0.0|"RT @kurteichenwald: @AchaPatricia You didnt read a lot of what I wrote pre-election, did you? Try these:https://t.co/JSN8Liptfchttps://t."
MattDocMartin|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
cowgirlup1a|qstafford50|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
cowgirlup1a|palmerreport|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
IapetusOrbit|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
janet_yackle|luvmom8702|0.0516|0.122|0.748|0.13|"RT @luvmom8702: @janet_yackle @TheCut President Obama and Hillary Clinton know, understand how wrong you&amp; trump are Women are strong in spi"
petersarsgaard|jonleeanderson|0.6808|0.145|0.578|0.277|RT @jonleeanderson: So the CIA says Kremlin hacked Hillary &amp; leaked intel to help Trump.He won &amp; will name a Putin friend Sec of State. Hav
ImForYOUAmerica|WayneDupreeShow|0.0|0.0|1.0|0.0|"RT @WayneDupreeShow: When Obama spoke with Russia in 2012, he said he would have leverage on hot mic, Hillary hit reset button with Putin.."
DoDFiredawg78|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
tigertrollz2|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
tigertrollz2||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
Kodie2038Donna|JKaetz|0.528|0.094|0.735|0.171|@JKaetz Bernie ALL TALK NO ACTION!!!!  WHY DIDNT HE STAND UP TO HILLARY AND THE DNC???  BECAUSE HE WAS PART OF THE GAME!  SMARTEN UP!
JuliaGhnaimat|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
ed_hooley|truthfeed|0.0|0.0|1.0|0.0|"British Diplomat ""I've Met The Wikileaks Informant and They're NOT Russian"" https://t.co/ocQMDX7il5 #ImWithHer #Hillary #maga"
Reinhard1934|LarryT1940|0.0|0.0|1.0|0.0|"RT @LarryT1940: Hey #Democrats, #Liberals, #MSM, #Hillary, #CIA &amp; #McCain, It wasn't #Russia. It was the message that blew #Hillary out of"
TerriGreenUSA|twitter|-0.0423|0.099|0.809|0.092|"We've already said no to #fakenews. DSW didn't deny anything wiki said, and there's still the investigation into Hi https://t.co/GMFsZntgHA"
ciji2016|charliekirk11|0.0|0.0|1.0|0.0|"RT @charliekirk11: Russia potentially being involved is a big deal, but where was the media when Hillary funded her entire staff with forei"
SawyerBrittain|gerfingerpoken|0.5696|0.0|0.735|0.265|RT @gerfingerpoken: (IBD) Why won't Hillary Get Prosecuted Like David Petraeus? - @IBDeditorials - #PJNET https://t.co/3lSPD7nnV2 - - https
SawyerBrittain|investors|0.5696|0.0|0.735|0.265|RT @gerfingerpoken: (IBD) Why won't Hillary Get Prosecuted Like David Petraeus? - @IBDeditorials - #PJNET https://t.co/3lSPD7nnV2 - - https
Duffy_1958|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
Duffy_1958|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
dougtgraham|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
dougtgraham||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
KevinMEaster|NakBananas|-0.2732|0.091|0.909|0.0|@NakBananas @YouTube there are different views on the subject. I still say Trump is unfit to be pres. Hillary's guilt doesn't change that.
DavidTravillia1|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
halfdollar54|YouTube|0.2577|0.0|0.865|0.135|HILLARY WONT EVEN HAVE MAJORITY OF VOTES ONCE THE DUST CLEARS https://t.co/9INvpMAXrZ via @YouTube
halfdollar54|youtube|0.2577|0.0|0.865|0.135|HILLARY WONT EVEN HAVE MAJORITY OF VOTES ONCE THE DUST CLEARS https://t.co/9INvpMAXrZ via @YouTube
LavaResistance|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
TeresaHutson1|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
TeresaHutson1|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
DAILYBLUEblog|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
sqhydusmhk3|sexdatehere2|-0.128|0.212|0.606|0.182|busty Hillary Scott lets her horny teacher fuck her sweet pussy https://t.co/7sOrV1jeBX
BJeanMohr1|twitter|0.507|0.122|0.612|0.266|"He's only good at insults, diplomacy is not his forte',HIllary is so much better at diplomacy. https://t.co/AjaSMhfQUE"
Me_iam_erica|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
sschrimp|corncob53|0.0|0.0|1.0|0.0|RT @corncob53: @LouDobbs @paulkrugman what's more de legitimizing than the Saudis $25 million contribution to HILLARY CLINTON? Krugman is a
PatHarr64573322|LovinPoulsbo|0.4019|0.094|0.749|0.157|RT @LovinPoulsbo: @HRCintheWild @katyperry  Love Hillary Clinton.  It won't be long before the entire US regrets not having her as our Pres
rickacoffman|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Gittoa1|youtube|0.0|0.0|1.0|0.0|Hillary calls for censorship https://t.co/Qv9C0Vklq1
Kdplayer13|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
jamie_roc|Ian56789|-0.4588|0.13|0.87|0.0|RT @Ian56789: Remember when Russian Hackers forced Hillary to wipe her server after being served with a Congressional Sub Poena to preserve
DoughnutJane|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
VikingsFan1964|billkooper|0.8126|0.0|0.697|0.303|@billkooper @GodH8sWindbags Obama won two consecutive terms. Hillary won with more than 2.5 million votes. The @ElectoralCollge hasn't voted
dssinojuli|ConstanceQueen8|0.7717|0.0|0.66|0.34|RT @ConstanceQueen8: Thank U 4 Sparing UsFrom Hillary Clinton Best Thanksgiving Ever Amen &amp; Amen #PresidentElectTrump #MA
AllWolvesMatter|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
BarrieNJ|IdiotDems|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
BarrieNJ|t|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
AnnTruwe|kylegriffin1|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
AnnTruwe|theatlantic|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
grammarox|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
DaleF3|eztempo|-0.7859|0.298|0.702|0.0|@eztempo @CNN Russia didn't do anything. Hillary's loss was her own damn fault. I'm not diving under my desk with my hands over my head.
nerfect|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
dawnsotolongo|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
dawnsotolongo|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
MelissaTT2000|LisaToddSutton|-0.3182|0.119|0.881|0.0|"@LisaToddSutton @KellyannePollsHillary say she lost, he is her president, willing to work w/ him. Get it yet, hon?https://t.co/i2gJFh3GUb"
MelissaTT2000|cnn|-0.3182|0.119|0.881|0.0|"@LisaToddSutton @KellyannePollsHillary say she lost, he is her president, willing to work w/ him. Get it yet, hon?https://t.co/i2gJFh3GUb"
LaurieRobert6|greggutfeld|0.0|0.0|1.0|0.0|"@greggutfeld @GregGutfeldShow Hillary dillary dock, her times run off the clock. Whitewater and email mishandled. Benghazi and foundation"
DAILYBLUEblog|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
Anfoooey|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
PatPatojson|FreedomChild3|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
PatPatojson|t|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
boris3324|davidfrum|0.0|0.0|1.0|0.0|"RT @davidfrum: Maybe it wasnt tactical, but I still dont understand why Hillary never said: Take off that pin, its not your flag, you P"
ZKondos|PatriotGeorgia|0.0|0.0|1.0|0.0|"@PatriotGeorgia @PatVPeters McCain, a Hillary/Obama/Soros surrogate must be removed from Chairman of the Armed Services committee"
riskmare|ezlusztig|0.0|0.0|1.0|0.0|RT @ezlusztig: From https://t.co/USXeAnLwWv
riskmare|theguardian|0.0|0.0|1.0|0.0|RT @ezlusztig: From https://t.co/USXeAnLwWv
PatDugan|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
MhMaximilian|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
MhMaximilian|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
titoriaanmol|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
conservogirl|RNRMississippi|-0.2263|0.215|0.642|0.143|"RT @RNRMississippi: Russians are Amazing: Set up a private server, rigged the primary, used BleachBit to violate a court order, then made"
amazinglyarden|twitter|-0.7626|0.267|0.733|0.0|HILLARY KNOWS SHIT YALL BUT NO WE NOW HAVE A CHEETO AS PRESIDENT WHO PROBABLY IS SECRETLY GAY WITH PUTIN https://t.co/KPYxj9ntdz
jwire|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
fakegreglambert|Eden_Eats|-0.5859|0.257|0.743|0.0|RT @Eden_Eats: Going on a hike without running into Hillary Clinton is bullshit.
edd79nyc|_CillaW|0.2732|0.0|0.92|0.08|RT @_CillaW: Agreed. It's all deep rooted sexism. Imagine if Hillary was elected &amp; doing half of the things Trump is right now. People woul
syl_pac|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/pyLGPjVyhG via @Change
syl_pac|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/pyLGPjVyhG via @Change
JohnVinhMiles|jackflackdaily|-0.4389|0.153|0.847|0.0|RT @jackflackdaily: Clinton Campaign Spent More Money Than Any Losing Campaign In US History!  https://t.co/QCwMkseXWc #Trump #makeamericag
JohnVinhMiles|redstate|-0.4389|0.153|0.847|0.0|RT @jackflackdaily: Clinton Campaign Spent More Money Than Any Losing Campaign In US History!  https://t.co/QCwMkseXWc #Trump #makeamericag
BizEnewsLive|Sterlingartz)hillary|0.4215|0.0|0.833|0.167|Retweeted Sterling J Sterling (@Sterlingartz):hillary clinton's lead in the popular vote swells to nearly 2.7... https://t.co/xEqDbVYxh8
BizEnewsLive|motherjones|0.4215|0.0|0.833|0.167|Retweeted Sterling J Sterling (@Sterlingartz):hillary clinton's lead in the popular vote swells to nearly 2.7... https://t.co/xEqDbVYxh8
tototch|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
FeistyTrumpette|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
lawnsports|benschwartzy|-0.5177|0.218|0.66|0.122|"RT @benschwartzy: It only took one FBI agent to ruin Nixon (Felt) and one to ruin Hillary (Comey). So, I'm very happy to see Trump making a"
aline260|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
aline260|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
tuckman_andrea|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
bloodinbritish3|Portosj81J|0.2263|0.0|0.924|0.076|RT @Portosj81J: If the CIA knew that Russia was behind hacking then why did Obama allow Hillary to use a private server with official secre
joneslisa|RamBoPirate|-0.4588|0.222|0.694|0.083|RT @RamBoPirate: Top 5 Reasons Hillary lost the Election:1-  She sux2-  She sux3-  She sux4-  She sux5-  She sux
Millenniumistic|freedemoparty|0.0|0.0|1.0|0.0|"RT @freedemoparty: PEOPLE'S LEADER MADAME PRESIDENT HILLARY CLINTON IS MARCHING TOWARDS ""THE WHITE HOUSE"" - Abdullah Al-Mahmud Jahangir htt"
PatriotRider|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
chris_jive|clwpaints|-0.4215|0.237|0.763|0.0|@clwpaints @MittRomney @joshromney    Do you think Hillary lies?  Just wondering
trishshirlaw|DineshDSouza|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
trishshirlaw|twitter|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
ScotiaMark|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
huffdini|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
LivingstonLD22|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
Sailfish157|Sherrishaw14|0.0|0.0|1.0|0.0|RT @Sherrishaw14: @whirrll @FredPecora @GOP @PatriotsOfMars @freep Hillary is the only one who can finish this https://t.co/uoRiqedjhA
Sailfish157|twitter|0.0|0.0|1.0|0.0|RT @Sherrishaw14: @whirrll @FredPecora @GOP @PatriotsOfMars @freep Hillary is the only one who can finish this https://t.co/uoRiqedjhA
paperrosie53|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
paperrosie53|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
Football__matri|blaubok|0.47|0.096|0.652|0.252|RT @blaubok: When her election was 98% certain - Hillary assured Trump - the election isn't riggedWhen she lost - the election was rigged
OldStudentnow|PBS|0.3481|0.047|0.85|0.103|@PBS @NewsHour How dare those Russian spread all that truth about #Hillary?  And why would they not want to deal with her corrupt legacy?
AgnesdeBerlimon|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
AgnesdeBerlimon|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
hillary_jar|JanethHdzSub|0.0|0.0|1.0|0.0|RT @JanethHdzSub: Cosas dificiles para harry: saludar y cantar al mismo tiempo#MTVStarsNiallHoran https://t.co/yL4f6ykE6D
hillary_jar|vine|0.0|0.0|1.0|0.0|RT @JanethHdzSub: Cosas dificiles para harry: saludar y cantar al mismo tiempo#MTVStarsNiallHoran https://t.co/yL4f6ykE6D
maryhowland7|WeNeedTrump|-0.802|0.31|0.69|0.0|@WeNeedTrump Hillary  made her  money from Morocco.Saudi. Bahrain.several  counties. She is mentally  ill from all her evil actions
Caranina01|Change|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/erYMV0p4oe via @Change
Caranina01|change|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/erYMV0p4oe via @Change
pambaker0208|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
caroljdavy|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
caroljdavy|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
macmcd|yourltldogtoo|0.0|0.0|1.0|0.0|RT @yourltldogtoo: .@amyklobuchar @washingtonpost Call on the #ElectoralCollege  to #DenyTrump and elect Hillary
hoseokway|maItinerecords|0.4019|0.0|0.838|0.162|RT @maItinerecords: hillary clinton flew all the way to hong kong to support twice https://t.co/Dsmufj6Xes
hoseokway|twitter|0.4019|0.0|0.838|0.162|RT @maItinerecords: hillary clinton flew all the way to hong kong to support twice https://t.co/Dsmufj6Xes
cakehler|swterry91|-0.4939|0.158|0.842|0.0|RT @swterry91: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money #tcot https://t.co/1b9uUjZ9lB
cakehler|dailycaller|-0.4939|0.158|0.842|0.0|RT @swterry91: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money #tcot https://t.co/1b9uUjZ9lB
marciebrowne|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
BizEctiveCTO|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
BizEctiveCTO|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
PrettySoftweb|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
PrettySoftweb|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
BizEnewsLive|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
BizEnewsLive|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
US_Conservatism|danbuter|-0.128|0.1|0.819|0.082|RT @danbuter: @nytimes @nytopinion Should do an article on the truth and lies of the New York Times. You'd get a whole series just on Hilla
dane0033|twitter|0.0|0.0|1.0|0.0|Or Hillary Clinton  https://t.co/JoiqJGM32e
ambinc1|umpire43|0.0|0.0|1.0|0.0|RT @umpire43: In Millwaukee day 5 of recount Hillary had 356000 votes thrown out for Fraud.Boxes in Millwaukee did not match poll books RUS
Newyorker2212|qstafford50|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
Newyorker2212|palmerreport|0.6249|0.0|0.746|0.254|"RT @qstafford50: Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,ta"
raklas|caveboyjones|0.5859|0.0|0.817|0.183|"@caveboyjones @infowars Actually, while MSM (FAKE NEWS) was predicting victory for Hillary, @infowars was accurately predicting Trump win."
suzost|pete03217|-0.8519|0.283|0.717|0.0|RT @pete03217: @lidiya_selwood @suzost @washingtonpost We see it but Dems choose not to see it. They are blind to all the horrible things H
Barbara4220|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
polyglotme|shayne571|-0.4767|0.14|0.86|0.0|@shayne571 @NoyzeSmythe @4everNeverTrump @caliwaterman @fawfulfan ur attack is same one Hillary used on Obama in 2008. it doesn't make sense
sherrysue66|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
sherrysue66|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
Michell8675309|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
mariemc11308417|IdiotDems|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
mariemc11308417|t|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
constantino_sam|pinterest|0.5423|0.163|0.485|0.352|I out of 3 Hillary supporters are  - ANTI HILLARY POLITICAL BUMPER FUNNY STICKER https://t.co/CcPjVHMd6h
sorceror43|andrea_manea|-0.4588|0.2|0.8|0.0|"@andrea_manea On Wall St, that was a Bernie issue.  Hillary wld have looked hypocritical."
forcerecon430|BrittPettibone|-0.8316|0.468|0.532|0.0|RT @BrittPettibone: Kellyanne Conway is battling a barrage of death threats from Hillary Supporters.#FridayFeelinghttps://t.co/0kLbme7ouQ
tony_c1967|thehill|-0.4767|0.181|0.819|0.0|"@thehill Worse than Hillary's? She made 33,000 emails go away w/ people pleading the 5th."
kitimi2|kitimi|-0.5267|0.207|0.793|0.0|Former U.S. Ambassador to Russia: Vladimir Putin Wanted Revenge on Hillary Clinton  Mediaite https://t.co/uTQJXE6evW
markguidry84|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
BrendaFiles2|umpire43|-0.5859|0.137|0.863|0.0|RT @umpire43: Hundreds of thousands of Fraud Hillary votes were foung in Detroit and in Millwaukee and in Philly. Did Russia do that to hel
stepvand|nytimesarts|0.3182|0.0|0.867|0.133|RT @nytimesarts: Madonnas speech about sexism put Hillary Clintons candidacy in fresh perspective. Discuss. https://t.co/uGEBHSXQOy https
stepvand|nytimes|0.3182|0.0|0.867|0.133|RT @nytimesarts: Madonnas speech about sexism put Hillary Clintons candidacy in fresh perspective. Discuss. https://t.co/uGEBHSXQOy https
JacksJungle|bfraser747|0.4215|0.0|0.865|0.135|"@bfraser747 if i were Putin, I'd think Hillary much easier to manipulate and control... Trump an unknown, America-first deal maker."
johnwalkergolf|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
conservogirl|manny_ottawa|-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
conservogirl||-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
SeattleHotDeals|seattleorganicrestaurants|0.0|0.0|1.0|0.0|RT #HighestRated most reliable business phone services: https://t.co/H35ipWVTWA and https://t.co/cdl60GAttE
JEKitten|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
JEKitten||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
starlady24|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
NJSappington|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: I repeat: I laid out what was going on with Russian campaign, based on leaks from European intel, before election: http"
Inductivist|washingtontimes|-0.8176|0.362|0.638|0.0|Hillary spends 2X as much as Trump ($1.2 b) &amp; lost miserably. Dems are terrible with money. https://t.co/Ozb7jQ72Q5
PeggyBurgess17|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
_antiheroine_|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
SiessChris|twitter|-0.7964|0.372|0.628|0.0|Nope. They were too busy making shit up to cover Hillary's fat ass. https://t.co/OevhAUkfbJ
bbeaty32|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
bbeaty32|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
SunnyAtTheGulf|RealMarkCole|0.0|0.0|1.0|0.0|RT @RealMarkCole: @brassmonkey3434 @peddoc63 did Russia put the earpiece in Hillary's ear or the teleprompter in her podium? https://t.co/L
SunnyAtTheGulf|luxmea|0.0|0.0|1.0|0.0|RT @RealMarkCole: @brassmonkey3434 @peddoc63 did Russia put the earpiece in Hillary's ear or the teleprompter in her podium? https://t.co/L
Bodisha|MichaelSollace|-0.9578|0.544|0.456|0.0|@MichaelSollace @ChrisCuomo awww... lol... poor lil fuck boy all sad there isn't gonna be a coronation for that evil bitch Hillary
ConservativeMag|conservativepapers|0.0|0.0|1.0|0.0|Heres What Could Happen if Hillary Clinton is Indicted or Steps Down https://t.co/eE4qxHNLIO #TeaParty #tcot
emiliocerejo|Quasar637|0.7363|0.0|0.735|0.265|"RT @Quasar637: @larryelder @EPS1991 don't forget she jailed Nakoula as part of the charade, Hillary &amp; Obama should both be jailed for that!"
TimKells1|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
ArtOfSamWood|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
GreenEyedLilo|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
mmedley41|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
HillaryBCrooked|VeteransTake|0.0|0.0|1.0|0.0|RT @VeteransTake: And Hillary said... #ArmyNavyGameDay #fakenews #MLSCup https://t.co/SZKW7OoHeB
HillaryBCrooked|twitter|0.0|0.0|1.0|0.0|RT @VeteransTake: And Hillary said... #ArmyNavyGameDay #fakenews #MLSCup https://t.co/SZKW7OoHeB
danbuter|nytimes|-0.128|0.107|0.805|0.088|@nytimes @nytopinion Should do an article on the truth and lies of the New York Times. You'd get a whole series just on Hillary.
ChefJennaMc|thehill|0.4382|0.0|0.822|0.178|"@thehill then you didn't pay attn to hillary's.She's been caught calling us deplorable,lying about emails is responsible for BENGAZI DEATHS!"
DeePSw31|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
PalinRevolution|SarahPalinUSA|0.0|0.0|1.0|0.0|RT @SarahPalinUSA: Rush reminds us ---&gt; https://t.co/VdGq41JjmZ https://t.co/BV9NwoEYvq
PalinRevolution|youngcons|0.0|0.0|1.0|0.0|RT @SarahPalinUSA: Rush reminds us ---&gt; https://t.co/VdGq41JjmZ https://t.co/BV9NwoEYvq
PoliticalPrick|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
PoliticalPrick|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
NonnieCon|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
seattle4events|seattleorganicrestaurants|0.0|0.0|1.0|0.0|RT #HighestRated most reliable business phone services: https://t.co/vmYdiP4phG and https://t.co/1V8TCObKNI
Genaritas1|Jason_Pollock|-0.1027|0.103|0.809|0.088|RT @Jason_Pollock: If you believed all the lies about Hillary then you played right into the hands of Russian hackers. Do you realize that
dms1013|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
vishnuduti|twitter|0.5927|0.0|0.845|0.155|"There had been a lot of foreign influence not only for Trump, but for Hillary, Quatar +Saudi Arabia are the good in https://t.co/eEYck73BaF"
Rickeyleetw|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
diewithbey|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
BloodyRed32|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
BloodyRed32||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
GrandCanyonPics|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
pie_jorge|intlspectator|0.8689|0.0|0.634|0.366|"RT @intlspectator: Hillary Clinton's popular vote lead now at 2.8 million votes, the greatest popular vote victory for presidential electio"
PaulieAbeles|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
PaulieAbeles|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
stickyfacts|youtube|0.0|0.0|1.0|0.0|Hillary Clinton Blew 1.2 Billion Dollars on Presidential Campaign!  https://t.co/JfiqvGdk3N
LKuehn4|summerbrennan|0.7003|0.0|0.707|0.293|"RT @summerbrennan: Joe Biden appealing to Trump voters. I wonder why? I hope good reasons, because https://t.co/1t6upiH0Tn https://t.co/Ypa"
LKuehn4|theatlantic|0.7003|0.0|0.707|0.293|"RT @summerbrennan: Joe Biden appealing to Trump voters. I wonder why? I hope good reasons, because https://t.co/1t6upiH0Tn https://t.co/Ypa"
LeslieNowicki1|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
NorbPeti|nytimes|0.3182|0.0|0.874|0.126|RT @nytimes: How a speech by Madonna about sexism put Hillary Clinton's candidacy in fresh perspective https://t.co/CqLswtts4u https://t.co
NorbPeti|nytimes|0.3182|0.0|0.874|0.126|RT @nytimes: How a speech by Madonna about sexism put Hillary Clinton's candidacy in fresh perspective https://t.co/CqLswtts4u https://t.co
conservogirl|PolitixGal|0.0|0.0|1.0|0.0|RT @PolitixGal: How Hillary really felt about the VOTERS! https://t.co/iPFPMyQcpk
conservogirl|twitter|0.0|0.0|1.0|0.0|RT @PolitixGal: How Hillary really felt about the VOTERS! https://t.co/iPFPMyQcpk
kailsss_10|sara_manbeck|0.0|0.0|1.0|0.0|"RT @sara_manbeck: ""What would you buy Hillary Clinton for Christmas?""-""Handcuffs"""
jacobspm|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
yourltldogtoo|amyklobuchar|0.0|0.0|1.0|0.0|.@amyklobuchar @washingtonpost Call on the #ElectoralCollege  to #DenyTrump and elect Hillary
cj_briomhar|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
lilradishn|twitter|-0.1935|0.259|0.547|0.194|"Nope! Hillary lost because if you are not a certifiable moron, she, of no personalty and/or clarity. She lost befor https://t.co/vNHkz3xG4M"
springerpappy|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
Debbie1228Hart1|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
safetyjedi|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
ColeHudson68|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
ColeHudson68|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
amerycarlson|asamjulian|-0.5267|0.201|0.738|0.061|"RT @asamjulian: It wasnt Russia, nor Comey. Hillary was an unlikable, uninspiring sociopath w/ no message and multiple legal problems. IT"
mgillaspie|corncob53|0.0|0.0|1.0|0.0|RT @corncob53: @LouDobbs @paulkrugman what's more de legitimizing than the Saudis $25 million contribution to HILLARY CLINTON? Krugman is a
BladeInTheHouse|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
Goodnightma|EcuadorDeb|0.0|0.0|1.0|0.0|"RT @EcuadorDeb: According to Podesta emails, her password was: Hillary.  My grandmother could hack that. Come on! https://t.co/uG1DmmlHdM"
Goodnightma|twitter|0.0|0.0|1.0|0.0|"RT @EcuadorDeb: According to Podesta emails, her password was: Hillary.  My grandmother could hack that. Come on! https://t.co/uG1DmmlHdM"
phil4gop|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
roqchrisy|DebAlwaystrump|0.5405|0.0|0.776|0.224|RT @DebAlwaystrump: HILLARY SELLS 20% OF USA URANIUM TO RUSSIAWHYDems must not be too worried about Russia sure Russia would want more
Queen_Raveen|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
KoolFreedom|SSReaney|0.0|0.0|1.0|0.0|"RT @SSReaney: @LMKay @bluepillXI @TheDemocrats ya know, I thought the exact same thing when Obama won...and we saw what he did; and Hillary"
trueiceman|WhosWyatt|0.5994|0.0|0.71|0.29|"@WhosWyatt @JohnUhan Trump supporter lol, and I'm assuming you voted for Hillary driving a Buick"
Marilunabeli|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
Marilunabeli|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
BarbaraLeeDeFra|change|0.0|0.0|1.0|0.0|THUS WE&gt;&gt;https://t.co/4gUj2vO5TO https://t.co/BehfHJqFt4
Betterw05759703|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: Think bout this: Allied intel servives investigating prez-elect 2 learn if he's Putin stooge in place 2 shatter NATO ht
roqchrisy|DebAlwaystrump|-0.5319|0.168|0.832|0.0|RT @DebAlwaystrump: RUSSIA HACKED CALIFORNIA 2GAVE THEM ALL DRIVERS LICENCES5.9 MILLION ILLEGALS LIVE IN SANCTUARY CITIES AND MADE T
popmuzikmofo|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
kaysunshine1252|CBSNews|0.4019|0.103|0.696|0.201|@CBSNews lol anyone or any country would favor Trump over Crooked Hillary. How many lies does Americans have to hear from her?OMG
washpress|nola|-0.7184|0.353|0.647|0.0|Hillary Clinton attacks 'fake news' in post-election appearance on Capitol Hill - https://t.co/uc3Ik4wESi https://t.co/MGHaD2aFJl
Awaken_the_46|FaceTheNation|0.0|0.0|1.0|0.0|@FaceTheNation @CarlaMoulton3 What's the endgame? Revote? Hillary/Pence? Any GOP is still a puppet &amp; Hillary will have endless clashes w/GOP
YourOpinionsAre|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
Anzers|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
jlpulice|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
jlpulice||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
MarthaLivingmar|mitchellvii|-0.1134|0.135|0.752|0.113|"@mitchellvii @DonWeldy And that is because the problems are never their fault, just ask Obama or Hillary."
cakehler|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
DrJADelgado|seanmdav|0.0|0.0|1.0|0.0|RT @seanmdav: And can you believe Putin made Hillary run more ads in Omaha than in Michigan and Wisconsin combined? Diabolical. https://t.c
DrJADelgado||0.0|0.0|1.0|0.0|RT @seanmdav: And can you believe Putin made Hillary run more ads in Omaha than in Michigan and Wisconsin combined? Diabolical. https://t.c
d_fucile|twitter|0.1511|0.111|0.756|0.133|"SHE NEEDS TO REALIZE SHE IS NOW JUST LIKE THE OTHERS IN THE PRIMARIES WHO ""LOST!""  HILLARY, YOU ARE A HASBEEN, A NO https://t.co/YtwW4cz6vg"
WayneABryant|umpire43|-0.4215|0.113|0.887|0.0|RT @umpire43: Before the SC shut down MI Recount. several hundred thousand Hillary votes disqualified as poll book and vote boxes did not m
diewithbey|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
JustineLee1993|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
JustineLee1993|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
roqchrisy|DebAlwaystrump|0.5405|0.0|0.776|0.224|RT @DebAlwaystrump: HILLARY SELLS 20% OF USA URANIUM TO RUSSIAWHYDems must not be too worried about Russia sure Russia would want more
kaiaka|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
MEDIATIONS99|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
WCurties|YouTube|-0.4278|0.215|0.673|0.112|Rush Limbaugh Plays Montage Of Hillary As A Purveyor Of FAKE NEWS https://t.co/pXTGWfL1yO via @YouTube
WCurties|youtube|-0.4278|0.215|0.673|0.112|Rush Limbaugh Plays Montage Of Hillary As A Purveyor Of FAKE NEWS https://t.co/pXTGWfL1yO via @YouTube
syqau|twitter|0.0|0.0|1.0|0.0|Hillary Clinton -- Russia Stole My Crown! ... https://t.co/H7oqYyiOSd
aaronhege|freddiedeboer|-0.4588|0.12|0.88|0.0|"RT @freddiedeboer: Russia forced Hillary's campaign to have one tenth as many canvassers in Michigan as John Kerry did 12 years earlier, cr"
beripsnicotti|LucidHuricane|-0.6792|0.411|0.589|0.0|RT @LucidHuricane: Whining Crying Rioting Hillary Millennial Theme Song!! https://t.co/wbLop5KvwL
beripsnicotti|twitter|-0.6792|0.411|0.589|0.0|RT @LucidHuricane: Whining Crying Rioting Hillary Millennial Theme Song!! https://t.co/wbLop5KvwL
The_Taxdude|johnnacalvillo|0.6908|0.0|0.695|0.305|"@johnnacalvillo @legendaryizaak Supporting crooked Hillary Clinton or socialist Bernie Sanders, favoring abortion and illegals amnesty."
mowser1970|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
xformed|gerfingerpoken|-0.34|0.179|0.714|0.107|RT @gerfingerpoken: (IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.
xformed|investors|-0.34|0.179|0.714|0.107|RT @gerfingerpoken: (IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.
g_rubylee2009|palmerreport|0.0|0.0|1.0|0.0|https://t.co/wozkylQANA
vatthepinters|daveweigel|-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
vatthepinters||-0.5719|0.239|0.667|0.094|"RT @daveweigel: ""Rejects politicization"" of intel, except when he calls for Hillary to be denied security briefings because email https://t"
caseywilder_|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
caseywilder_||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
pearlygates101|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
yceek|yceek|0.0|0.0|1.0|0.0|RT @yceek: Farewell --- Hillary Clinton  - LAST Big Rally https://t.co/5RzMP0IlOj
yceek|twitter|0.0|0.0|1.0|0.0|RT @yceek: Farewell --- Hillary Clinton  - LAST Big Rally https://t.co/5RzMP0IlOj
texliberty|facebook|0.0516|0.124|0.702|0.174|I've concluded that if Hillary Clinton attacked Satan there are a good number of people on the right who would... https://t.co/VPTMJjMouz
suzost|RealMarkCole|0.3111|0.166|0.628|0.206|@RealMarkCole MSM &amp; Dems don't know how to handle Trump! Fake News! Alt RT! Comey Russia Yes it was definitely Russia! No it's Hillary! 
rickydiva227|nytimes|0.3182|0.0|0.874|0.126|RT @nytimes: How a speech by Madonna about sexism put Hillary Clinton's candidacy in fresh perspective https://t.co/CqLswtts4u https://t.co
rickydiva227|nytimes|0.3182|0.0|0.874|0.126|RT @nytimes: How a speech by Madonna about sexism put Hillary Clinton's candidacy in fresh perspective https://t.co/CqLswtts4u https://t.co
apple_butter|parisswade|0.4153|0.137|0.664|0.199|RT @parisswade: WOW TREY GOWDY HAS HIT A TIME BOMB HERE WITH HILLARY AND HER HENCHMEN !!KEEP AT IT TREY GOWDY !!!https://t.co/bvgmk9iqqK
apple_butter|usapoliticstoday|0.4153|0.137|0.664|0.199|RT @parisswade: WOW TREY GOWDY HAS HIT A TIME BOMB HERE WITH HILLARY AND HER HENCHMEN !!KEEP AT IT TREY GOWDY !!!https://t.co/bvgmk9iqqK
jen_thorson|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
lightlady|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
NicolasRobidoux|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
ThorntonScout|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
Marmel|TheBaxterBean|-0.3182|0.113|0.887|0.0|"RT @TheBaxterBean: REMINDER: Hillary Clinton lost Michigan by only 10,704 votes. Detroit has 513,000 registered voters &amp; turnout declined ("
Brendybob|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
echogaffney|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/Gtc7J2OSli
connieSuver|CarmineZozzora|-0.3007|0.254|0.594|0.152|"RT @CarmineZozzora: Hillary's criminal activity on her unsecured server putting America's national security at risk wasn't a problem, but D"
Angie_B2011|7b00f339f69e48f|0.0|0.0|1.0|0.0|"RT @7b00f339f69e48f: @TuckerCarlson @realDonaldTrump @FoxNews offered 5 cents on a dollar for Hillary's fireworks!!! ""I thought I""de get a"
9951jackson|BigDuhie1955|0.0|0.0|1.0|0.0|@BigDuhie1955 obama now joined in on the hacking order Cia to look in to the hacking.hillary should be session first thing he does
glover53a|youtube|-0.34|0.255|0.745|0.0|Hillary Clinton to Face A Firing Squad-FBI director https://t.co/NCtgWwlSHk
JagbusAnne|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
JagbusAnne|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
kldreams61|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
msjbe20a|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
jvargasnow|PeakOfTruth|0.25|0.124|0.677|0.199|RT @PeakOfTruth: Anyone who honestly believes Russia is responsible for #Hillary getting rolled is 2 dumb to continue to draw oxygen https:
bigdaddydoggie|MeghanMG|-0.6124|0.208|0.792|0.0|@MeghanMG @MightyChin @Tablavi @keksalamander And CROOKED Hillary lost to him. I guess its not  saying much about her to lose to a nunce.
bwtanker|GabbyInCa|0.0|0.0|1.0|0.0|"@GabbyInCa @SpecialKMB1969 @60Minutes @netanyahu @realDonaldTrump  unlike Obama &amp; Hillary, told the press things tht should never been said"
rigormortis1961|JudgeJeanine|0.5927|0.0|0.845|0.155|@JudgeJeanine Hillary deserves a bag of coal for Christmas but that's even too good for her so I'd give her just the bag. 
artandmusicmom|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/rEFrGwb2xZ via @Change
artandmusicmom|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/rEFrGwb2xZ via @Change
Redskins_4me|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
katemccloudsays|wolfgangfaustX|-0.6904|0.263|0.737|0.0|"@wolfgangfaustX @JohnMerlyn618 @dave_cpt @Stevenwhirsch99  Intel comm. not trust Hillary? HA,HA. Now they have POTUS who doesn't trust them!"
Hillary_Rdz|valtrevy|0.0|0.0|1.0|0.0|@valtrevy rale ya te extrao 
gregfahlgren|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
StopHillary01|dailycaller|-0.6705|0.314|0.686|0.0|Morning Joe' Calls Out Hillary For 'Fake News' Warning | The Daily Caller https://t.co/ymw30lESuP #politics
LifeWinnersOnly|dailycaller|-0.6124|0.313|0.688|0.0|Hillary Campaign Ignored Staffer Who Predicted She'd Lose | The Daily Caller https://t.co/VEWulSEspS #breaking
ConservNationA|dailycaller|-0.6705|0.314|0.686|0.0|Morning Joe' Calls Out Hillary For 'Fake News' Warning | The Daily Caller https://t.co/Vz2iixsLRd #politics
patriotnewsone|foxnews|0.0|0.0|1.0|0.0|What's next for Hillary? Latest moves indicate Clinton won't fade away |  #breaking  https://t.co/bys9QI8zHw
Trillion3|CNN|0.0|0.0|1.0|0.0|@CNN https://t.co/kRF9EM73lH https://t.co/C4iFdwmehA
Trillion3|thegatewaypundit|0.0|0.0|1.0|0.0|@CNN https://t.co/kRF9EM73lH https://t.co/C4iFdwmehA
kenene1|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
KCDurling|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Bluebugaboo2|twitter|0.0|0.0|1.0|0.0|You didn't  get it Hillary sold our uranium illegally toPutin without consulting congress. That's a crimenot conf https://t.co/52ObDB3rhW
GreerSusan|change|0.0|0.0|1.0|0.0|Federal Registrar of the U.S. Electoral College: Did you know that there is still a way to elect Hillary Clinton... https://t.co/lkLwsgmSoG
mimi_x4|TheTobster111|0.7717|0.0|0.712|0.288|"RT @TheTobster111: Legal precedence says that you don't hold new elections, the results of old are overturned. Add to that winning popular"
fixedopsjack|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
fixedopsjack|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
carlaho15238423|realjunsonchan|0.4076|0.133|0.632|0.235|"RT @realjunsonchan: -@KellyannePolls completely rekts Rotten Hillary. Lol. This is how America should be governed, spend less, win more. Ni"
EventosJlcervys|Change_Mex|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/09juKINLoN va @Change_Mex
EventosJlcervys|change|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/09juKINLoN va @Change_Mex
CaptainM72|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
CaptainM72|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
SGTROCKUSMC82|twitter|-0.3182|0.161|0.839|0.0|Why didn't they figure this out before the election that Hillary lost? https://t.co/mwxPUkHahn
dkcollins27|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
JarrettOSmith|canjcat|0.7804|0.0|0.771|0.229|@canjcat @Reince That's why WE call you liberated. YOU believe what you hear instead of what you know. Hillary won the election says MSM. HA
jmingerson725|HillaryClinton|-0.6908|0.26|0.65|0.09|@HillaryClinton @timkaine @billclinton @ChelseaClinton HILLARY I urge you to stand up and fight like hell for your rightful seat in the WH
connieSuver|CarmineZozzora|-0.2991|0.15|0.791|0.058|RT @CarmineZozzora: They didn't care about Hillary's unsecured server of classified and top secret info in her backyard - but who dared to
geh4osu|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
gomi0526|soledadobrien|0.0|0.0|1.0|0.0|@soledadobrien @TrinityNYC @dmitryzaksAFP @HillaryClinton Hillary was born a decade or so too early.
maryjamesblige|twitter|0.0|0.0|1.0|0.0|Hillary said this in every debate but woah buddy those emails https://t.co/gyI0ojcuZT
JoshuaMPatton|latest_com|-0.6115|0.222|0.778|0.0|RT @latest_com: Harvard Study: Hillary Clinton Received The Most Negative Coverage in 2016Campaign https://t.co/M8munNI1xo https://t.co/Ug
JoshuaMPatton|latest|-0.6115|0.222|0.778|0.0|RT @latest_com: Harvard Study: Hillary Clinton Received The Most Negative Coverage in 2016Campaign https://t.co/M8munNI1xo https://t.co/Ug
kee_raje|KjThaMonarch|0.0|0.0|1.0|0.0|RT @KjThaMonarch: How imma be When they announce trump for president #election2016 #trumptrain #hillary #comedy #jokes https://t.co/fGWIGg
kee_raje|t|0.0|0.0|1.0|0.0|RT @KjThaMonarch: How imma be When they announce trump for president #election2016 #trumptrain #hillary #comedy #jokes https://t.co/fGWIGg
jtrevizo1013|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
devinedianakins|GodandtheBear|0.2584|0.0|0.912|0.088|RT @GodandtheBear: I'm not crazy about Hillary is an understatement as to what I feel towards that psychopath. Him being one doesn't change
AllWolvesMatter|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
thatgirlsandra5|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
TheSoniaV|OccupyDemocrats|0.128|0.0|0.914|0.086|RT @OccupyDemocrats: #Breaking News: Russian Hacks Just Gave Courts Legal Precedent To Replace Trump With Hillary https://t.co/SqdHfv4GYo
TheSoniaV|occupydemocrats|0.128|0.0|0.914|0.086|RT @OccupyDemocrats: #Breaking News: Russian Hacks Just Gave Courts Legal Precedent To Replace Trump With Hillary https://t.co/SqdHfv4GYo
Alllwftopic|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
CobyRayan|VeronicaGriman|-0.5319|0.177|0.823|0.0|RT @VeronicaGriman: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/aaWkrfbssx https://t.co/XghezX5He8
CobyRayan|truthfeed|-0.5319|0.177|0.823|0.0|RT @VeronicaGriman: This Video Details How Hillary Blew $1.2 BILLION to LOSE the White House https://t.co/aaWkrfbssx https://t.co/XghezX5He8
stilllwithher|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
constantino_sam|pinterest|-0.5319|0.378|0.428|0.194|HILLARY FOR PRISON 2016 - ANTI HILLARY POLITICAL BUMPER FUNNY STICKER https://t.co/RTgtHPXzCt
ka4_trump|Republiicunts|0.0772|0.122|0.741|0.138|@Republiicunts @kristinw2is @RealNathanHale @mitchellvii @NateSilver538 Hillary lost the Electoral College. It's time to accept the result
Mr_Liva|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
glover53a|youtube|-0.6369|0.426|0.574|0.0|'Hillary Clinton exposed for the death of thousands.' https://t.co/cvky5aAYTO
lwestsd|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
peacelovedixie|DPRK_News|0.6705|0.113|0.604|0.283|RT @DPRK_News: Supreme Leader Kim Jong-Un telegrams congratulations to Russian president Vladimir Putin on defeat of venomous fish-wife Hil
emccoy_writer|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
oldcrookedhouse|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
amandaspleas|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
EducWoman|charliekirk11|-0.5719|0.201|0.727|0.073|"RT @charliekirk11: Hillary blames ""fake news"" for her lossFunny, the media is the only reason clinton did as well as she did,  She would"
cala_1111|truthfeed|-0.4069|0.163|0.837|0.0|Did #RussianHackers HIDE the State of Wisconsin from Hillary Clinton? Social Media Chimes in! https://t.co/Ka10yoNRlF
richard19079|2ALAW|0.0|0.0|1.0|0.0|RT @2ALAW: The American Nightmare Coming To An End  01/20/17#Trump#Hillary https://t.co/vh7ngOZxWX
richard19079|twitter|0.0|0.0|1.0|0.0|RT @2ALAW: The American Nightmare Coming To An End  01/20/17#Trump#Hillary https://t.co/vh7ngOZxWX
rachyohreally|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
JETMEDIA2|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
c5wired97|umpire43|-0.4215|0.113|0.887|0.0|RT @umpire43: Before the SC shut down MI Recount. several hundred thousand Hillary votes disqualified as poll book and vote boxes did not m
MariusLecter|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
BTW_LOL|gerfingerpoken|-0.34|0.179|0.714|0.107|RT @gerfingerpoken: (IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.
BTW_LOL||-0.34|0.179|0.714|0.107|RT @gerfingerpoken: (IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.
BugsbJr|PrisonPlanet|-0.7845|0.317|0.683|0.0|"RT @PrisonPlanet: Ed Klein: Hillary cried inconsolably, blamed Comey &amp; Obama for not doing enough to stop FBI investigation. https://t.co/K"
BugsbJr|t|-0.7845|0.317|0.683|0.0|"RT @PrisonPlanet: Ed Klein: Hillary cried inconsolably, blamed Comey &amp; Obama for not doing enough to stop FBI investigation. https://t.co/K"
Noahsbet|charliekirk11|-0.5106|0.13|0.87|0.0|RT @charliekirk11: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
MRSTXFabFace|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
kimberlymontse1|standupgyrl|0.0|0.0|1.0|0.0|@standupgyrl @TravisRuger as if Hillary's choices would be any different #HelloOligarchy
Apatriot11|softwarnet|-0.2732|0.091|0.909|0.0|"RT @softwarnet: ""FBI and CIA""Podesta was warned in 2008 to use encryption, Hillary didn't, DNC didn't, Obama's OPM didn't - those who igno"
Hispanics16|usapoliticstoday|-0.6221|0.316|0.684|0.0|Forget Russia! Reince Priebus Just Pointed Out Why Hillary Really Lost! https://t.co/Xt9RsXNLZY https://t.co/uxa0pvcUAc
jakesCove_US|Flirman1983|-0.8402|0.321|0.679|0.0|"RT @Flirman1983: @JohnKStahlUSA They lied, cheated and stoled the Dem. nomination and have the audacity to say Fake News caused Hillary' lo"
pammcbide55|DebAlwaystrump|0.5405|0.0|0.776|0.224|RT @DebAlwaystrump: HILLARY SELLS 20% OF USA URANIUM TO RUSSIAWHYDems must not be too worried about Russia sure Russia would want more
swaglee214|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
nicks847|dick_nixon|0.0|0.0|1.0|0.0|RT @dick_nixon: I got called an asshole when I wrote this. https://t.co/5GZYN5250r
nicks847|thedailybeast|0.0|0.0|1.0|0.0|RT @dick_nixon: I got called an asshole when I wrote this. https://t.co/5GZYN5250r
coreyhaines|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
honorverity|ragdog1|-0.6679|0.233|0.767|0.0|RT @ragdog1: @Khanoisseur Hillary told Americans! They did not listen! Now you fools we pay the price. Loosing our country!
latest_com|latest|-0.6115|0.25|0.75|0.0|Harvard Study: Hillary Clinton Received The Most Negative Coverage in 2016Campaign https://t.co/M8munNI1xo https://t.co/Ugc1pi6xkW
WhosWyatt|trueiceman|-0.8271|0.372|0.628|0.0|.@trueiceman @JohnUhan because my b u ick would look fuckin sick faggot you probably voted for Hillary
WakeUpCanada1|ed_hooley|-0.7269|0.337|0.663|0.0|RT @ed_hooley: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/RKOyB0S2vR
WakeUpCanada1|nytimes|-0.7269|0.337|0.663|0.0|RT @ed_hooley: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/RKOyB0S2vR
rockrexx|NorthFalcon74|-0.4019|0.114|0.886|0.0|RT @NorthFalcon74: @Portosj81J @Dewblue1 Notice nobody is saying *what* was hacked. The fact is it was Hillary Clinton's server. End of sto
wtf_imtooold|MJB_SF|0.0|0.0|1.0|0.0|RT @MJB_SF: and that is: Elect Hillary Clinton. #AuditTheVote #hamiltonelectors https://t.co/2Rke9GAdRY
wtf_imtooold|twitter|0.0|0.0|1.0|0.0|RT @MJB_SF: and that is: Elect Hillary Clinton. #AuditTheVote #hamiltonelectors https://t.co/2Rke9GAdRY
CarlNyberg312|ggreenwald|-0.5362|0.154|0.846|0.0|On what issue did GOP attack Hillary Clinton as too far to the Left? When did she take these positions?@ggreenwald
edmecka|edmecka|-0.6124|0.357|0.643|0.0|Hillary Campaign Ignored Staffer Who Predicted Shed Lose |  https://t.co/59ja18sKiG via @edmecka
edmecka|dailycaller|-0.6124|0.357|0.643|0.0|Hillary Campaign Ignored Staffer Who Predicted Shed Lose |  https://t.co/59ja18sKiG via @edmecka
springerpappy|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
TuxiTix4|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
cb55uic|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
volpappaw|DailyCaller|-0.8126|0.359|0.641|0.0|RT @DailyCaller: Shooting The Wrong Messenger  Morning Joe Calls Out Hillary Clinton For Hiding Behind Fake News https://t.co/gq71mB
volpappaw|t|-0.8126|0.359|0.641|0.0|RT @DailyCaller: Shooting The Wrong Messenger  Morning Joe Calls Out Hillary Clinton For Hiding Behind Fake News https://t.co/gq71mB
mtighe15|MrDane1982|0.1007|0.161|0.714|0.125|"RT @MrDane1982: 40 yrs of fighting for us, this time we fight for her until she have enough ground to stand on! The best thing Hillary can"
frostdeeds|Seriousman67|0.4019|0.0|0.828|0.172|RT @Seriousman67: @bessbell @realDonaldTrump Hillary has had saudi support and massive donations from them
BugsbJr|DebAlwaystrump|0.5405|0.0|0.776|0.224|RT @DebAlwaystrump: HILLARY SELLS 20% OF USA URANIUM TO RUSSIAWHYDems must not be too worried about Russia sure Russia would want more
LoveMyRedCat|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/p4zEjyg3Ro via @Change
LoveMyRedCat|linkis|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/p4zEjyg3Ro via @Change
close_jonathan|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
starry_galaxies|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
MsLiveat5|Justin_CMeck|0.2732|0.0|0.913|0.087|@Justin_CMeck @CNN well I did hear an analyst on PBS both Hillary Clinton and Donald Trump had a office in the same building N/ Delaware
realrobottrump|vox|-0.2023|0.114|0.815|0.071|By how it feels I want to cut and run in Libya and #iraq leaving our country  https://t.co/CenZD1I7XO
ka3byz|umpire43|-0.5859|0.147|0.853|0.0|RT @umpire43: When it is now proven fact and on record that thousands of Fraud Hillary votes in 3 recount states lets INVESTIGATE THAT
Hillary_Rdz|valtrevy|0.0|0.0|1.0|0.0|RT @valtrevy: @Hillary_Rdz JAJAJAJA maldita desesperada ya casi me voy para all
Hnurse07|LindaSuhler|0.4404|0.0|0.847|0.153|RT @LindaSuhler: A good time to mention Hillary Clinton's REAL link to Russia...#RussianHackingShe transferred our uranium to Putin...FOR
petersonaj|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
SaysSheToday|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
shannoncaraker|twitter|0.0|0.0|1.0|0.0|Hillary be like.....#Trump2016 #RussiaHacking #RedNationRising https://t.co/7jMKm1ESmP
YoYoDietByBy|AlessaAndreadis|0.7322|0.0|0.722|0.278|"RT @AlessaAndreadis: @LouDobbs @realDonaldTrump has a charm about him that so many Americans enjoy, something Hillary lacked entirely. (But"
TINKLEY1|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
staggerlee420|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
frostdeeds|BentleyforTrump|-0.2893|0.204|0.651|0.145|RT @BentleyforTrump: @bessbell @realDonaldTrump A 1000 Times better than fucking Crooked ass Hillary! #QueenOfTheLies and #QueenOfTheFlies
ImmoralReport|dreamedofdust|0.4574|0.0|0.85|0.15|RT @dreamedofdust: #HillaryForPrison ! https://t.co/OWXj4jLsry They started with me in the 1990s then. (If you're convinced that Hillary is
ImmoralReport|reddit|0.4574|0.0|0.85|0.15|RT @dreamedofdust: #HillaryForPrison ! https://t.co/OWXj4jLsry They started with me in the 1990s then. (If you're convinced that Hillary is
Word_Made_Death|gerfingerpoken2|-0.5106|0.18|0.82|0.0|RT @gerfingerpoken2: #Benghazi Mom Patricia Smith Targets Serial Liar Hillary https://t.co/KVO6ImiEzS - American Thinker - #PJNET 999 - htt
Word_Made_Death|americanthinker|-0.5106|0.18|0.82|0.0|RT @gerfingerpoken2: #Benghazi Mom Patricia Smith Targets Serial Liar Hillary https://t.co/KVO6ImiEzS - American Thinker - #PJNET 999 - htt
Animal1984Farm|DRUDGE_REPORT|-0.8137|0.277|0.723|0.0|@DRUDGE_REPORT Obamas hate the Clintons they don't want them near in WH. DNC hacks only made Hillary &amp; her inner circle look bad not obama
Chericrane11|marlins360|0.3612|0.148|0.604|0.248|@marlins360 @tonyposnanski @JoelNihlean @realDonaldTrump No actually Hillary won the most votes
doogsadavis|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
2eyesnears|cristinalaila1|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
2eyesnears|twitter|-0.3182|0.247|0.753|0.0|RT @cristinalaila1: Hillary Clinton lost again #TriggeredIn4Words https://t.co/zgXW7Yt5Ty
espresso_4|"washingtonpost,"|0.4019|0.0|0.87|0.13|"@washingtonpost, hopefully, at the same time, they'll investigate the extent and consequences of the hacking of Hillary's email server."
Wayne5Juan|DiAlegna|0.0|0.0|1.0|0.0|RT @DiAlegna: #ImStillNotOver Hillary saying things she doesn't actually mean. #NeverHillary ';&gt; https://t.co/0PCzV6wTpD
Wayne5Juan|twitter|0.0|0.0|1.0|0.0|RT @DiAlegna: #ImStillNotOver Hillary saying things she doesn't actually mean. #NeverHillary ';&gt; https://t.co/0PCzV6wTpD
Humanbeingish|jfgroves|0.25|0.073|0.813|0.114|"RT @jfgroves: Wait, the woman who offered blowjobs to vote for Hillary is complaining about sexism in the music industry? Lol. https://t."
Humanbeingish||0.25|0.073|0.813|0.114|"RT @jfgroves: Wait, the woman who offered blowjobs to vote for Hillary is complaining about sexism in the music industry? Lol. https://t."
Travii_Johnson|Change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/eZH4N1CQUd via @Change
Travii_Johnson|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/eZH4N1CQUd via @Change
Espen414|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
pjwilb|PhxKen|0.0|0.0|1.0|0.0|RT @PhxKen: HILLARY CLINTON SAYS WE HAVE TO MANY GUNS IN AMERICA. I SAY WE HAVE TO MANY CLINTONS. https://t.co/Bvmbz6uHiN
pjwilb|twitter|0.0|0.0|1.0|0.0|RT @PhxKen: HILLARY CLINTON SAYS WE HAVE TO MANY GUNS IN AMERICA. I SAY WE HAVE TO MANY CLINTONS. https://t.co/Bvmbz6uHiN
ReelTPJ|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
opticspolitics|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
opticspolitics|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
safeminefield|Im_ConnorKelley|0.7901|0.0|0.696|0.304|"@Im_ConnorKelley @realDonaldTrump @NBCNightlyNews @CNN ""Hillary won by 2.83 million *FAKE* votes"". There fixed it for you. You're welcome!"
ShirlZitting|LisaToddSutton|-0.4767|0.154|0.846|0.0|@LisaToddSutton @Deplorable_B @Battlep431 @KellyannePolls Hack this hack that. Poor Hillary was hacking out a cough every word she spoke.
texascornhuske1|PiceaLives|0.8126|0.0|0.641|0.359|"@PiceaLives @blakehounshell @politico Spruceass is the kind who supports corruption and lawlessness, like Hillary and Obama. Scum liberal."
ellenichen|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
polyglotme|shayne571|0.3612|0.0|0.894|0.106|"@shayne571 Bernie led progressive consensus, wasn't part of establishment like Hillary was, so it was naturally harder for him to pass laws."
Confederate265|ReversingASD|0.0|0.0|1.0|0.0|RT @ReversingASD: Fox News LiveHILLARY BELONGS IN JAIL! TREY GOWDY VS HILLARY CLINTON US News Today https://t.co/tuqjfyKmNF via @youtube
Confederate265|youtube|0.0|0.0|1.0|0.0|RT @ReversingASD: Fox News LiveHILLARY BELONGS IN JAIL! TREY GOWDY VS HILLARY CLINTON US News Today https://t.co/tuqjfyKmNF via @youtube
rockrexx|Portosj81J|0.2263|0.0|0.924|0.076|RT @Portosj81J: If the CIA knew that Russia was behind hacking then why did Obama allow Hillary to use a private server with official secre
susanmanners|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Luchadora213|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
hii1701|TrinityNYC|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
hii1701|t|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
4freedomamerica|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
MI2CA2|peddoc63|0.1531|0.084|0.812|0.104|RT @peddoc63: Do you care that Hillary sold 20% of our Uranium to Russians? Or that Obama lied to pass Iran Deal &amp; Obamacare &amp;that he paid
SusanCarver19|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
tonic516|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
MrPhotoDave2k|mikandynothem|0.7324|0.0|0.755|0.245|"RT @mikandynothem: So far, the ""recount"" isn't going so well for Hillary. Trump GAINS votes in Wisconsin! #TrumpCabinetBand #MAGA #tcot ht"
GretchenInOK|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Bry574|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
Bry574|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
PaulieAbeles|charliekirk11|-0.5106|0.13|0.87|0.0|RT @charliekirk11: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
steveg1425|Pappiness|0.5859|0.0|0.833|0.167|"RT @Pappiness: Just a subtle reminder that if #RussianHackers helped Hillary win, The GOP Oversight Committee would investigate her for tre"
melwusa|brunelldonald|-0.6486|0.29|0.627|0.082|@brunelldonald Only if Hillary Clinton is rightfully Charged with the same and many other Felony Charges as well at https://t.co/FJaSnALEAT
melwusa|twitter|-0.6486|0.29|0.627|0.082|@brunelldonald Only if Hillary Clinton is rightfully Charged with the same and many other Felony Charges as well at https://t.co/FJaSnALEAT
DonnaRo86165010|RepStevenSmith|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
DonnaRo86165010|dailycaller|-0.4939|0.167|0.833|0.0|RT @RepStevenSmith: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/Y6BazF4OsJ v
Chambord22|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
curtvendel|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
blessedone333|iparker6642|-0.5255|0.166|0.834|0.0|@iparker6642 @atticalocke @Vote4TrumpPrez she voted for the traitor Hillary who's treatment of poor black Haitians is LEGENDARY! #FullMoron
RebeccaKovalich|DailyMail|-0.6542|0.328|0.672|0.0|RT @DailyMail: Hillary's policy director warned her she could lose election 'but everyone ignored him' https://t.co/AcRG3xTO8r
RebeccaKovalich|dailymail|-0.6542|0.328|0.672|0.0|RT @DailyMail: Hillary's policy director warned her she could lose election 'but everyone ignored him' https://t.co/AcRG3xTO8r
JBax52|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
JBax52|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
AtsukoNatsume|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
AtsukoNatsume|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
luvruthy|ArianeBellamar|0.0|0.0|1.0|0.0|RT @ArianeBellamar:  b4 Partisan! Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/CMOS
luvruthy|t|0.0|0.0|1.0|0.0|RT @ArianeBellamar:  b4 Partisan! Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/CMOS
Yosbones|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
Luchadora213|LindaSuhler|0.4404|0.0|0.847|0.153|RT @LindaSuhler: A good time to mention Hillary Clinton's REAL link to Russia...#RussianHackingShe transferred our uranium to Putin...FOR
TheRick35|bfraser747|-0.6901|0.222|0.778|0.0|"RT @bfraser747:  ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."" ~ @GovMikeHu"
bridget4kicks|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
mmsahaj|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
mmsahaj|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
glenda045|bennydiego|0.2382|0.0|0.911|0.089|RT @bennydiego: It's funny how Hillary's private server was such a major issue but President-elect talking to world leaders on his private
blackandgold43|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
stateroute1776|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
TCCKatherine1|change|0.0|0.0|1.0|0.0|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/zsRXJt9dgW
DEALMEEIN2016|MarcosBreton|0.178|0.138|0.703|0.159|"RT @MarcosBreton: If it was the same ""old"" news, but with Hillary Clinton as the winner, YOU and every Repbulican would be SCREAMING for an"
katgrneyes|charliekirk11|-0.5106|0.13|0.87|0.0|RT @charliekirk11: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
tomotb|America_1st_|-0.6901|0.222|0.778|0.0|"RT @America_1st_: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candi"
Patrioticgirl86|2ALAW|-0.3182|0.223|0.777|0.0|RT @2ALAW: @LeahR77 @SenJohnMcCain @LindseyGrahamSC Hillary Sees A Ghost https://t.co/EOvIdoE4iU
Patrioticgirl86|twitter|-0.3182|0.223|0.777|0.0|RT @2ALAW: @LeahR77 @SenJohnMcCain @LindseyGrahamSC Hillary Sees A Ghost https://t.co/EOvIdoE4iU
akhsilom|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
nolbol|S1776frdm|-0.9186|0.519|0.417|0.064|"RT @S1776frdm: Hillary Sucked at everything except Treason Corruption Pay4PlayKindness of Spirit Racism, Hate 4 Average Citizens--https:/"
nolbol||-0.9186|0.519|0.417|0.064|"RT @S1776frdm: Hillary Sucked at everything except Treason Corruption Pay4PlayKindness of Spirit Racism, Hate 4 Average Citizens--https:/"
4gatoscuba|DLasAmericas|0.0|0.0|1.0|0.0|@DLasAmericas @realDonaldTrump Y siguen en el negocio? Esa encuestadora dijo que hillary ganaba elecciones con 41% y Trump perdia con 37%.
NatlTimes|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
Frances_davis1|TheMarkRomano|0.0|0.0|1.0|0.0|"RT @TheMarkRomano: Hey Hillary, just an FYI...Letting 30-year-old Pajama Boy @RobbyMook run your Presidential campaign, was not such a gr"
gerfingerpoken|IBDeditorials|-0.34|0.199|0.682|0.119|(IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.co/kNFLEno9Tb
gerfingerpoken|investors|-0.34|0.199|0.682|0.119|(IBD) If Hillary Signed Form OF-109 she committed Felony - @IBDeditorials #PJNET 999 https://t.co/127jNePgDg https://t.co/kNFLEno9Tb
Ivorysnow3567|DineshDSouza|-0.1943|0.216|0.671|0.113|@DineshDSouza @HillarysAmerica No idea why people refused to SEE TRUTH. I worked hard for trump  if Hillary we&gt; be Islam Nation peeps sleep
Shari_Cookson|ShepsMom|0.8122|0.135|0.509|0.356|"RT @ShepsMom: Hillary lost by a questionable 80k votes, won 3 Million more popular votes, yet #Trump still claims big win as excuse for #ru"
Anonymouthpiece|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
Anonymouthpiece|t|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
BarbaraLeeDeFra|Change&gt;&gt;SIGN|0.4981|0.0|0.832|0.168|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/zcpgCCW5gt via @Change&gt;&gt;SIGN &amp; SHARE
BarbaraLeeDeFra|change|0.4981|0.0|0.832|0.168|Electoral College: Make Hillary Clinton President on December 19 - Sign the Petition! https://t.co/zcpgCCW5gt via @Change&gt;&gt;SIGN &amp; SHARE
TischaSingh|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
TischaSingh|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
Trinidadiyon|twitter|-0.5829|0.166|0.834|0.0|"America has the most backward ass democracy, if you know Russia influenced a whole election why not do a revote? Hi https://t.co/4N7Lz7Js8k"
MaryTrinetti|occupydemocrats|0.128|0.0|0.889|0.111|Russian Hacks Just Gave Courts Legal Precedent To Replace Trump With Hillary - https://t.co/ZjKCPyYBRK
sheri_scary|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
Jonathan_Estes|Domm_G_|0.5859|0.0|0.817|0.183|@Domm_G_ inside climate control vs outside in the elements... you must've also knew Hillary was going to win
blueskymountain|bennydiego|0.2382|0.0|0.911|0.089|RT @bennydiego: It's funny how Hillary's private server was such a major issue but President-elect talking to world leaders on his private
gerfingerpoken|t|0.0|0.0|1.0|0.0|Enabler Hillarys Actions Speak Louder Than Trumps Words - Flopping Aces - https://t.co/zGKDjKzaBM-  https://t.co/Sl1y6adA8U #MAGA
JB__Cali|thegatewaypundit|-0.4939|0.151|0.849|0.0|Sen. D'Amato Drops Bomb: Hillary Allowed Russia to Take Ownership of US Uranium to Sell to Iran (Video) https://t.co/XgK0rpS5Ia
LindaHenrichsen|discus74|-0.3818|0.126|0.874|0.0|RT @discus74: @AlisonSpalding2 @SharNeal Hillary and Bill have manipulated our Gov't to feed their ostentatious lifestyles and become power
Hispanics16|usapoliticstoday|-0.4767|0.193|0.807|0.0|"Joe Scarborough: HILLARY CLINTON COST HILLARY CLINTON THE ELECTION, Not Fake News https://t.co/vaw8FwlP1r https://t.co/jgIBtonzJa"
JaniceTXBlessed|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
KevinAParker1|VeteransTake|0.0|0.0|1.0|0.0|RT @VeteransTake: And Hillary said... #ArmyNavyGameDay #fakenews #MLSCup https://t.co/SZKW7OoHeB
KevinAParker1|twitter|0.0|0.0|1.0|0.0|RT @VeteransTake: And Hillary said... #ArmyNavyGameDay #fakenews #MLSCup https://t.co/SZKW7OoHeB
brandon120|twitter|-0.1531|0.108|0.811|0.081|We need to admit that Bernie Sanders was right and should be president now.  Hillary was a mistake of a candidate. https://t.co/WoXcWmFoS5
perry46_Shirley|PaulKinkel|-0.101|0.111|0.796|0.093|RT @PaulKinkel: Hillary sets up a homebrew server with less security than I have in my home Dems complain about #RussianHackers. Yup.
debdasp|charliekirk11|-0.765|0.369|0.631|0.0|@charliekirk11 @wendyvoss media will lose money..hillary alrleady lost a billion and Clinton fdn is losing money too
HeykbBennett|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
LMCraig|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
m_q_d_|VABVOX|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
m_q_d_|t|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
LKinTX|ETGilmour|-0.0258|0.226|0.599|0.175|@ETGilmour @GtaThoughts @HeyTammyBruce EVERYONE thought Hillary would win incl Putin. Russians hacked to undermine Hillary's presidency
ghw91|VABVOX|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
ghw91|t|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
SpringsRaff|Einsteinrevisit|-0.5994|0.205|0.795|0.0|RT @Einsteinrevisit: @dcexaminer  When the @FBI  was asked if Russia had hacked Clinton Server...Team Hillary and MSM SHOUTED no proof. Yet
PupTart|mmpadellan|0.0|0.0|1.0|0.0|RT @mmpadellan: Think about it.Ever see a 70yr old man UNHINGED 2 the point of grade-school taunts?Hillary CALLED it on #RussianHackers.
ClaydYila|JohnWascavage|0.0|0.0|1.0|0.0|"RT @JohnWascavage: Do you ever imagine that every morning Hillary Clinton wakes up and goes out into a field and sings ""Rose's Turn"" to Ame"
hbbtruth|carinabergfeldt|-0.3818|0.14|0.86|0.0|@carinabergfeldt MT @nypost - #Hillary campaign spent twice as much as #Trump on her losing presidential campaign. https://t.co/TKYcPLKovq
hbbtruth|twitter|-0.3818|0.14|0.86|0.0|@carinabergfeldt MT @nypost - #Hillary campaign spent twice as much as #Trump on her losing presidential campaign. https://t.co/TKYcPLKovq
DarinDorsey4|mitchellvii|-0.5905|0.211|0.714|0.076|@mitchellvii @ZarkoElDiablo @HillaryClinton I rarely disagree will @mitchellvii but the problem with Hillary was she was Hillary Clinton!!!
MizCoretta|AdamsFlaFan|-0.3612|0.167|0.739|0.094|"RT @AdamsFlaFan: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/wokIcX3tph via @crooksandliars"
MizCoretta|crooksandliars|-0.3612|0.167|0.739|0.094|"RT @AdamsFlaFan: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/wokIcX3tph via @crooksandliars"
paolo_sf|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
paolo_sf|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
JackGattanella|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
ClaydYila|rolandscahill|-0.3346|0.16|0.694|0.146|RT @rolandscahill: I think we all need a cathartic 11 o'clock number by Hillary Clinton to help get through this insanity. A Rose's Turn fo
mabian|HumanistReport|-0.4019|0.31|0.69|0.0|RT @HumanistReport: Why did Hillary Clinton lose?
connocrat|lukeoneil47|-0.6597|0.293|0.707|0.0|RT @lukeoneil47: The Democrats hacked the election and emails ...but to make Hillary lose https://t.co/QstENq3dbl
connocrat|twitter|-0.6597|0.293|0.707|0.0|RT @lukeoneil47: The Democrats hacked the election and emails ...but to make Hillary lose https://t.co/QstENq3dbl
AFRICANAMERICA1|KailiJoy)Hillary|0.7003|0.095|0.603|0.302|Retweeted Kaili Joy Gray (@KailiJoy):Hillary Clinton's under no obligation to save us. She tried. And we... https://t.co/N6MsjX4mrF
AFRICANAMERICA1|facebook|0.7003|0.095|0.603|0.302|Retweeted Kaili Joy Gray (@KailiJoy):Hillary Clinton's under no obligation to save us. She tried. And we... https://t.co/N6MsjX4mrF
PatPatojson|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
HShadeeth|Fiolanastacia|-0.296|0.155|0.845|0.0|"@Fiolanastacia Hillary, y no sigo viva y perreando Jajajajajaja me quede dormida como 5 minutos ajaja"
DragonTat2|TheXclass|-0.1139|0.126|0.874|0.0|RT @TheXclass: @SierraCynic @KatyGerhold @BLUpfront @popsknox @SenSanders They don't want a revote. They want Hillary to ascend to the thro
Bronxgirl418|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
jeweltyme|gerfingerpoken2|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
jeweltyme|floppingaces|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
kellyfirehorse|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
roqchrisy|spacedrogue|-0.4215|0.157|0.843|0.0|RT @spacedrogue: #Assange addresses the lies spread by #Hillary months before the election:https://t.co/pd69uOW8YqRussia hack is #FakeNew
roqchrisy|t|-0.4215|0.157|0.843|0.0|RT @spacedrogue: #Assange addresses the lies spread by #Hillary months before the election:https://t.co/pd69uOW8YqRussia hack is #FakeNew
mimi_x4|MelindaThinker|0.2023|0.0|0.833|0.167|RT @MelindaThinker: Russian interference with the election could give courts legal authority to install Hillary https://t.co/By58AeeOe3
mimi_x4|huffingtonpost|0.2023|0.0|0.833|0.167|RT @MelindaThinker: Russian interference with the election could give courts legal authority to install Hillary https://t.co/By58AeeOe3
qstafford50|palmerreport|0.7163|0.0|0.728|0.272|"Prominent attorney sues FBI for improperly favoring Donald Trump over Hillary Clinton https://t.co/m2cwaX2p00 the fight,take it to SCOTUS!!!"
Lynnsmith63Lynn|twitter|-0.4019|0.184|0.816|0.0|Holy SH*T BALLS. NSA Hacked DNC&amp;HILLARY JUDGE NAPOLITANO WAS INFORMED BY NSA https://t.co/ErUXacA4KC
Pauldias73|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
AFRICANAMERICA1|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
aliezirasch1|RealMarkCole|0.0|0.0|1.0|0.0|RT @RealMarkCole: @brassmonkey3434 @peddoc63 did Russia put the earpiece in Hillary's ear or the teleprompter in her podium? https://t.co/L
aliezirasch1|luxmea|0.0|0.0|1.0|0.0|RT @RealMarkCole: @brassmonkey3434 @peddoc63 did Russia put the earpiece in Hillary's ear or the teleprompter in her podium? https://t.co/L
mdsmelser|538politics|-0.6808|0.259|0.741|0.0|RT @538politics: Hillary Clinton's weakness in the Midwest is really the Democratic Party's weakness in the Midwest. https://t.co/gdAdESwM9
mdsmelser|t|-0.6808|0.259|0.741|0.0|RT @538politics: Hillary Clinton's weakness in the Midwest is really the Democratic Party's weakness in the Midwest. https://t.co/gdAdESwM9
baileelee|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
SilkWithDiamond|JudicialWatch|0.0|0.0|1.0|0.0|RT @JudicialWatch: In this country our leaders are bound by the rule of law. Hillary Clinton must be held accountable for her actions.http
MelonieFerry|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
Lee_in_Iowa|SwissTriple_M|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
Lee_in_Iowa|palmerreport|0.0|0.0|1.0|0.0|"RT @SwissTriple_M: @socialcivility @posybass1 https://t.co/P2y62B8SmT 70% voted early in FLA, more D than R, early exit P showed 1/2"
muttsandersbro|kurteichenwald|0.0|0.0|1.0|0.0|"@kurteichenwald @ericgarland ""But Hillary!"""
GrumpyOldSport|FiveThirtyEight|0.5719|0.1|0.68|0.22|"According to Yahoo, I'm 80% favorite to win my playoff game. About where @FiveThirtyEight had Hillary near end of Oct. What could go wrong?"
johnykakes|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
johnykakes||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
Smize21|realDonaldTrump|-0.5439|0.164|0.836|0.0|RT @realDonaldTrump: Hillary said she was under sniper fire (while surrounded by USSS.) Turned out to be a total lie. She is not fit to lea
abbaeema41|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""It was PresidentObama, along with Hillary Clinton, that came up with the 'Russian reset button"" ~ @AllenWest#JudgeJeani"
LeftAmerican|MMFlint|-0.6966|0.2|0.8|0.0|RT @MMFlint: Have you heard a ONE Dem leader scream about this? Imagine if Cuba hacked in to throw the election to Hillary? What would Repu
FMixmaster|charliekirk11|-0.5106|0.13|0.87|0.0|RT @charliekirk11: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
cussetabraswell|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
ksc12991|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
ksc12991||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
scott_stalker2|AmericanMex067|-0.6486|0.22|0.735|0.045|"RT @AmericanMex067: She had fake news backing her, DOJ, Obama - spent $1.2 billion &amp; still lost. Russia had nothing 2 do w/it.https://t.co"
Revolution41157|GodandtheBear|-0.8225|0.388|0.612|0.0|"RT @GodandtheBear: Hillary is the worst of bad people, a wolf in sheep's clothing. https://t.co/wy3ux6sLx9"
Revolution41157|twitter|-0.8225|0.388|0.612|0.0|"RT @GodandtheBear: Hillary is the worst of bad people, a wolf in sheep's clothing. https://t.co/wy3ux6sLx9"
zztopf450|immigrant4trump|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
zztopf450|twitter|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
DellaMelton57|twitter|0.2263|0.0|0.917|0.083|"Nothing surprises me about Obama &amp; his henchmen. Thru Hillary, he thought he'd be getting a 3rd term to put his las https://t.co/QCx1Ewfu9J"
cesario_brenden|MatthewOhman|0.0|0.0|1.0|0.0|@MatthewOhman Hillary is that you 
carolyn_pearl|Ian56789|-0.4588|0.13|0.87|0.0|RT @Ian56789: Remember when Russian Hackers forced Hillary to wipe her server after being served with a Congressional Sub Poena to preserve
JeffreyGuterman|MJBodary|-0.8687|0.471|0.529|0.0|"RT @MJBodary: You are disgusting human waste, JefferyGuterman.Hillary Clinton is a liar and a crook!#shameful https://t.co/g9zzvEYhMp"
JeffreyGuterman|twitter|-0.8687|0.471|0.529|0.0|"RT @MJBodary: You are disgusting human waste, JefferyGuterman.Hillary Clinton is a liar and a crook!#shameful https://t.co/g9zzvEYhMp"
susancrawshaw|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
susancrawshaw||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
TruthEqualsFact|GOP|0.0|0.0|1.0|0.0|"The @GOP in the Electoral College must cast their votes to Hillary Clinton, America's REAL PRESIDENT. https://t.co/ntx2A3AoKT"
TruthEqualsFact|twitter|0.0|0.0|1.0|0.0|"The @GOP in the Electoral College must cast their votes to Hillary Clinton, America's REAL PRESIDENT. https://t.co/ntx2A3AoKT"
southparkzombie|m|0.0|0.0|1.0|0.0|https://t.co/SZOxrBgEkq
braden_rose|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
ghostknife78|pudcast245|-0.6486|0.185|0.815|0.0|"@pudcast245 @SaintsTailgate @vivelafra I bet u Trump hacks who blieve Hillary is a killer 4real, also believe Batman is based on real events"
truther_dare|TimRunsHisMouth|0.6654|0.0|0.729|0.271|@TimRunsHisMouth @Cernovich did Hillary win? Why are you still using her to deflect?!
jtrevizo1013|KailiJoy|-0.6331|0.283|0.609|0.108|RT @KailiJoy: Hillary Clinton's under no obligation to save us. She tried. And we screamed EMAILS!!!!!! and complained that she's just not
Patrioticgirl86|LeahR77|-0.5106|0.163|0.837|0.0|RT @LeahR77: Tweedle Dee &amp; Tweedle Dumb @SenJohnMcCain  &amp; @LindseyGrahamSC Should Be Investigating Hillary's Home Brewed Server #FakeNews #
springerpappy|PeakOfTruth|0.25|0.124|0.677|0.199|RT @PeakOfTruth: Anyone who honestly believes Russia is responsible for #Hillary getting rolled is 2 dumb to continue to draw oxygen https:
theaterboy520|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
ed_hooley|nytimes|-0.7269|0.379|0.621|0.0|Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/RKOyB0S2vR
MissCrawford88|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
MsRachelWolf|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
jllundqu|Lynn_Rose1|0.0|0.0|1.0|0.0|@Lynn_Rose1 @ba613 @SammyHains tell that to Hillary. She exploded Libya and the state dept is largely cover for CIA ops in those lands.
b_drone|correctthemedia|-0.296|0.136|0.864|0.0|RT @correctthemedia: Hillary wants us to stop paying attention to news about child trafficking. https://t.co/KYy3bQLd5X
b_drone|twitter|-0.296|0.136|0.864|0.0|RT @correctthemedia: Hillary wants us to stop paying attention to news about child trafficking. https://t.co/KYy3bQLd5X
tkdnaz5|nia4_trump|-0.7096|0.258|0.742|0.0|RT @nia4_trump: Hillary blames Russia &amp; #FakeNews for her lossReality Check it was the Scandals Corruption Collusion &amp; Divisivenesshttps:
5Against1Eight3|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
5Against1Eight3||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
scott_stalker2|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
MayerDmayer6940|veggie64_leslie|-0.5574|0.204|0.796|0.0|RT @veggie64_leslie: A delusional story about why Hillary lost that captures the lack of responsibility of Clinton and her followers  http
amnesty11|gerfingerpoken2|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
amnesty11|floppingaces|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
beth_deitchman|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
dr_ashok_m|twitter|-0.1531|0.114|0.795|0.091|"But is has to be #Russia that got Donna Brazille to cheat for #Hillary in debates, she is such an innocent buffalo, https://t.co/R6WXDOkuHA"
gamecocksSecE|heyjoshhaines|-0.3595|0.122|0.878|0.0|".@heyjoshhaines paid protestors? I'm speaking of Hillary, Podesta, DNC colluding to disrupt election against Bernie try and keep up!"
Gan1Nancy|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
Gan1Nancy|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
lanasunb|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
emmandaluz|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
emmandaluz|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
TriCrescent|DaysOfTrump|-0.5994|0.196|0.804|0.0|"RT @DaysOfTrump: #AmericaFirst Patriots inside USgov are waging a civil war w international socialists (Hillary, Soros..) that have infiltr"
Michelem1998|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
logophobe|ByYourLogic|-0.4847|0.125|0.875|0.0|RT @ByYourLogic: i still don't understand why hillary clinton didn't go super saiyan. i'm 60 years old and make six figures to write about
ValerieEllenLe1|kurteichenwald|-0.2382|0.22|0.67|0.11|"RT @kurteichenwald: No offense, @chucktodd, but when u say no one was sure Russia behind hack pre-election, shows u need to read more. http"
TheMuseCompels|JYSexton|0.0|0.0|1.0|0.0|RT @JYSexton: This isn't about Donald Trump or Hillary Clinton. It's about sovereignty. It's about rights.
Margag_|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
consmover|DrMartyFox|-0.2732|0.123|0.877|0.0|RT @DrMartyFox: IF #RussianHackers Helped #Trump They Did By Exposing What The #DishonestMedia Was ConcealingCorrupt #Hillaryhttps:
FatherShaggy|late2game|-0.296|0.095|0.905|0.0|@late2game I thought there was a threshold of implausibility for that. Running in the woods: no pic. Running into Hillary in the woods: pic.
2eyesnears|lionelverney|0.0|0.0|1.0|0.0|RT @lionelverney: Wait ~ what ~ Hillary is a woman ? Chelsea Handler urges women to unite: 'Let's open our arms to each other'https
MstrWaterbender|HumanistReport|-0.4019|0.124|0.876|0.0|RT @HumanistReport: The left will never learn their lesson because they're still scrambling to find a scapegoat for Hillary Clinton's terri
meemo51956|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
tpuskas98|LibertyLivesHer|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
tpuskas98|vivaliberty|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
debyoungblood|drturpin|0.7351|0.0|0.721|0.279|RT @drturpin: Retweeted I'm still w/Hillary (@Mon9lem):That's wonderful news. Scott Dworkin thank you for not allowing these... https://t
debyoungblood||0.7351|0.0|0.721|0.279|RT @drturpin: Retweeted I'm still w/Hillary (@Mon9lem):That's wonderful news. Scott Dworkin thank you for not allowing these... https://t
brittreneehall|AdamParkhomenko|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
brittreneehall|nydailynews|0.0|0.0|1.0|0.0|RT @AdamParkhomenko: Hillary Clinton sent a thank-you note to a 103-year-old Long Island woman who voted for her https://t.co/3pRFSF3goq ht
trumptup2016|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
sleeper9|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
Kmich718|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
Kmich718|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
Ramo_Jr|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
JeremyHimli|shoahnuffin1|-0.4639|0.223|0.666|0.111|@shoahnuffin1 Just yesterday Trump laughed when the crowd chanted about jailing Hillary and said we don't care about that anymore. Sucker.
Col_Connaughton|youtube|0.0|0.0|1.0|0.0|Hillary Clinton is Deteriorating AGAIN! https://t.co/EUS46dseOo #hillary #clinton #degenerate #downhill
JanFrye|worldnetdaily|-0.2263|0.174|0.826|0.0|Hillary pleads to dismiss lawsuit against her https://t.co/beq2kJnkGv via @worldnetdaily
JanFrye|wnd|-0.2263|0.174|0.826|0.0|Hillary pleads to dismiss lawsuit against her https://t.co/beq2kJnkGv via @worldnetdaily
winstar1k|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
OteroReog51|iorch_athosfcab|0.0|0.0|1.0|0.0|"RT @iorch_athosfcab: @CNNEE pero los Wikileaks dijeron cosas ciertas acerca de Hillary, la Cia siempre busca crear caos."
constantino_sam|pinterest|-0.4648|0.216|0.784|0.0|Give Hillary's Dad a Condom - ANTI HILLARY PRO TRUMP POLITICAL BUMPER STICKER https://t.co/arlCLdvLSt
MarshaMc1203|Molloromma|0.6369|0.101|0.614|0.285|@Molloromma Hillary won by over 2 1/2 million votes. Trump is a minority president. He lost the popular vote.
frenchiesrock|hale_razor|-0.6925|0.206|0.794|0.0|"RT @hale_razor: Every U.S poll had Hillary crushing Trump in Wisconsin, but Putin's ground game in Madison knew it was close so he hacked p"
j_breents|SheWhoVotes|-0.7096|0.211|0.789|0.0|"RT @SheWhoVotes: If Hillary was complicit in Russian treason the way Donald is, I'd rightly turn on her. This should be unacceptable to *al"
JohnEhmet|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
Demontialto|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
conservogirl|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
conservogirl|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
wes332012|TheMichaelRock|-0.2732|0.208|0.679|0.113|RT @TheMichaelRock: My 8yo just kicked my ass in Battleship. This must be what Hillary Clinton feels like.
MariaClass|change|0.0|0.0|1.0|0.0|"Over 4.8 million people have signed the petition ""Electoral College: Make Hillary Clinton President"". https://t.co/y9xppRaMZF"
wy8162|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
wy8162|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
TheAuraWah|Vickigr81567276|0.0|0.0|1.0|0.0|@Vickigr81567276 @healRonaldTrump @FoxNews who can get a boner for Hillary? Not even all the world's Viagra can do that.
PatPatojson|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
ChrisLanzetti|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
georgeshannon11|JudgeJeanine|-0.4707|0.226|0.668|0.106|@JudgeJeanine i still cannot believe people are so stupid  about hillary Yes it was hard for me to spell that name
Eazy_Arts|VABVOX|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
Eazy_Arts|t|0.6908|0.0|0.778|0.222|"RT @VABVOX: 8) Hillary Clinton's popular vote lead (2,835,808) is now FIVE TIMES larger than Al Gore's was in 2000 (543,895): https://t.co/"
heywealtright|PrisonPlanet|-0.3527|0.202|0.665|0.133|@PrisonPlanet Lol Hillary's gonna get her Russian War one way or another huh? What's Mensch's salary?
arawis|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: The Democrats all debate who's going to get out of Hillary's way first, except for VERMONT'S OWN BERNIE SANDERS, who...get"
PoliticalMinion|MittRomney|0.6908|0.0|0.725|0.275|Hillary save America from Trump release your electors to vote 4 a normal Republican like @MittRomney https://t.co/1QIJU04q5b via @HuffPost
PoliticalMinion|huffingtonpost|0.6908|0.0|0.725|0.275|Hillary save America from Trump release your electors to vote 4 a normal Republican like @MittRomney https://t.co/1QIJU04q5b via @HuffPost
BarrieNJ|twitter|0.6322|0.0|0.771|0.229|The Nate Silver that predicted Hillary would win in a monumental landslide?  That Nate Silver? https://t.co/nUaXgBN3aB
kevpand|twitter|0.128|0.088|0.805|0.107|"For the Hillary fans, here are some nice scenic views from a county she lost to Bernie in the primaries and then to https://t.co/PJ7PU4K9Pa"
TrumpDyke|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
Wyohawk|immigrant4trump|-0.9136|0.432|0.568|0.0|"RT @immigrant4trump: Hillary ""Liar of the Year""  Blames Fake News, and Russia for Lost, Electoral Landslide Loss to Trump 308 VS 232 #mag"
jauremom|brandongroeny|-0.5106|0.13|0.87|0.0|RT @brandongroeny: Where was media outcry when Hillary sold out US for millions from foreign donors to the Clinton Foundation? That is fo
BryonnyMackay|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
BryonnyMackay|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
Evasabe|stylistkavin|-0.7269|0.289|0.711|0.0|RT @stylistkavin: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/pqjurgsNw7 #SistersinArms @Madonna @Hillar
Evasabe|nytimes|-0.7269|0.289|0.711|0.0|RT @stylistkavin: Madonna and Hillary: Witch and Nasty Woman as Sisters in Arms https://t.co/pqjurgsNw7 #SistersinArms @Madonna @Hillar
DuplexHaver|AliAbunimah|-0.3265|0.171|0.727|0.102|"RT @AliAbunimah: .@JoyAnnReid before and after Hillary, due to Democrat incompetence not Pootin, lost election. https://t.co/89GH9UWVdA"
DuplexHaver|twitter|-0.3265|0.171|0.727|0.102|"RT @AliAbunimah: .@JoyAnnReid before and after Hillary, due to Democrat incompetence not Pootin, lost election. https://t.co/89GH9UWVdA"
chuckc247|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
gcofmt42|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
RobertSAdcock|WeNeedTrump|-0.296|0.091|0.909|0.0|"RT @WeNeedTrump: Liberals crack me up when they call Trump ""Putin's puppet"" with no evidence. Yet millions of dollars donated to Hillary is"
PatPatojson|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: Hillary's secret $2.35M Russian Connection was so crooked, even the #CorruptMedia had to covered it. #UraniumOnehttps://t."
RamonleeRoush1|JudgeJeanine|0.3639|0.191|0.571|0.239|@JudgeJeanine  you think you're so funny wisecracking on Hillary Clinton what have you done that makes you so special I think you're STUPID!
ArgotMay|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
kingtynk|DineshDSouza|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
kingtynk|twitter|-0.3182|0.173|0.827|0.0|RT @DineshDSouza: The reason Hillary lost is not Russia--it's this guy https://t.co/tERRJGv05E
WileyCoyote9999|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
robdobber81|NBCNews|0.0|0.0|1.0|0.0|"@NBCNews Unlike Bill and Hillary, new cabinet members likely produced something rather than taking cash from foreign countries."
ChrisRocca2|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
RonTamber|gerfingerpoken2|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
RonTamber|floppingaces|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
gigi2my4|LVNancy|0.5719|0.0|0.791|0.209|"RT @LVNancy: #RussianHackers IF sore-Loser, Hillary had won, would we be having this conversation?#SundayMorning #TRUMP#AmericaFirst"
zwwwara|GeorgeTakei|0.5719|0.0|0.875|0.125|"RT @GeorgeTakei: If the CIA had found Russia had helped Hillary, and she had won by a razor thin margin, how do you suppose the GOP and its"
DuplexHaver|MaxBlumenthal|0.0|0.0|1.0|0.0|RT @MaxBlumenthal: .@AliAbunimah @JoyAnnReid What we've learned here is that Putin took out Hillary but Hillary did not take out Qaddafi. h
tadpoledrain|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
bikerbd|immigrant4trump|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
bikerbd|twitter|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
lorilpeabody|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
NadeemFayad|pmaft|-0.7351|0.292|0.708|0.0|RT @pmaft: If You Applied Hillary Clintons Logic On The Real Victims Of War ToRape https://t.co/ONxNk1b6aw https://t.co/EftLaJifhX
NadeemFayad|antifeministtech|-0.7351|0.292|0.708|0.0|RT @pmaft: If You Applied Hillary Clintons Logic On The Real Victims Of War ToRape https://t.co/ONxNk1b6aw https://t.co/EftLaJifhX
Redskins_4me|syqau|-0.5106|0.292|0.708|0.0|"RT @syqau: Rotten Sicko Hillary Clinton's ""fact checkers""... https://t.co/HQrGztLSiA"
Redskins_4me|twitter|-0.5106|0.292|0.708|0.0|"RT @syqau: Rotten Sicko Hillary Clinton's ""fact checkers""... https://t.co/HQrGztLSiA"
valtrevy|Hillary_Rdz|0.0|0.0|1.0|0.0|@Hillary_Rdz JAJAJAJA maldita desesperada ya casi me voy para all
nicegirlnks|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
MichaelDeitz1|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
MichaelDeitz1||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
trubdub88|BetteMidler|0.4201|0.0|0.883|0.117|"RT @BetteMidler: Donald Trump calls on Hillary to shut down her foundation. Meanwhile, were all still begging him to choose a more natural"
ArtPar17|hrtablaze|-0.644|0.226|0.774|0.0|RT @hrtablaze: Remember when wikileaks revealed that Primaries were rigged for Hillary? Are the Russians to blame for that too?https://t
ArtPar17||-0.644|0.226|0.774|0.0|RT @hrtablaze: Remember when wikileaks revealed that Primaries were rigged for Hillary? Are the Russians to blame for that too?https://t
BoatBonnie|vivelafra|-0.4019|0.241|0.623|0.136|RT @vivelafra: MEET THE AMATEUR: @ChuckTodd's buffoonish loyalty to #Hillary is beyond embarrassing &amp; destroys the credibility of @MeetTheP
1isten_up|PaulKinkel|-0.101|0.111|0.796|0.093|RT @PaulKinkel: Hillary sets up a homebrew server with less security than I have in my home Dems complain about #RussianHackers. Yup.
LavaResistance|nia4_trump|0.0|0.0|1.0|0.0|"RT @nia4_trump: #PodestaEmails more proof of Hillary's Russian Connections. ""Grassley Letter"" to Loretta Lynch. #CorruptMedia let this stor"
xraysoheil|WordSmithGuy|-0.743|0.24|0.76|0.0|RT @WordSmithGuy: Hillary Clinton spent twice as much as Trump in losing presidential bid. Negative TV ads don't connect with people. https
Freedom55555553|Justin_CMeck|0.0516|0.223|0.581|0.197|"@Justin_CMeck @CNN No, unfortunately it was lost when the bathroom server was moved. We just have to trust Hillary and Bill.. bless them"
ladieann|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
hillary_bentley|twitter|0.0|0.0|1.0|0.0|089#___#____#__#__#__ https://t.co/H86sVBsLDE
TroyCoby|TroyCoby|0.0|0.0|1.0|0.0|RT @TroyCoby: Hillary Clinton has been drinking a lot... https://t.co/vPJh1ZkOFN
TroyCoby|twitter|0.0|0.0|1.0|0.0|RT @TroyCoby: Hillary Clinton has been drinking a lot... https://t.co/vPJh1ZkOFN
jessicat_f|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
Twisty58|America_1st_|-0.6901|0.222|0.778|0.0|"RT @America_1st_: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candi"
JkbComic|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
akborough|conservativetribune|0.0772|0.0|0.894|0.106|Hillary Won&amp;#8217;t Even Have Majority of Votes Once the Dust Clears https://t.co/vonygLWGMx
2006ta|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
TheRick35|immigrant4trump|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
TheRick35|twitter|-0.7269|0.253|0.747|0.0|RT @immigrant4trump: Hillary Loser of the Year  The first woman to lose the same election twice #maga #trump #maga https://t.co/bzjEk58v7R
PatPatojson|jimlibertarian|0.4939|0.0|0.856|0.144|"RT @jimlibertarian: Donald Trump only works 4 we the people and America,Hillary Clinton on the other hand is a Chinese/Russian agent,she so"
NoMediaSpin|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
2dsnarow|Deeliberatrix|0.1779|0.16|0.642|0.198|@Deeliberatrix @LisaToddSutton @KellyannePolls electoral map proves won by a landslide get over it. Hillary sucked
PaulieAbeles|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
TheOxyCon|seanmdav|0.5267|0.085|0.704|0.211|"RT @seanmdav: So Russia is the reason Hillary ""You're Likable Enough"" Clinton lost in 2008? That seems like pretty big news. https://t.co/L"
TheOxyCon|luxmea|0.5267|0.085|0.704|0.211|"RT @seanmdav: So Russia is the reason Hillary ""You're Likable Enough"" Clinton lost in 2008? That seems like pretty big news. https://t.co/L"
FKWONdane|TrinityNYC|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
FKWONdane|t|0.0|0.0|1.0|0.0|RT @TrinityNYC: https://t.co/FE3kumenP9CNN
GaryfRiera|JohnLeguizamo|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
GaryfRiera|t|0.0|0.0|1.0|0.0|RT @JohnLeguizamo: Over 4 million have already asked the electoral college to elect @HillaryClinton as president on Dec 19. https://t.co/gh
txconservgirl|twitter|0.5423|0.0|0.632|0.368|Another article praising HillaryLibs never learn#wakeuplibs https://t.co/18KQTcTcQ8
JReiter18|JohnEkdahl|0.0|0.0|1.0|0.0|RT @JohnEkdahl: Hillary leaves her server open to hacking. Obama rolls over on his belly for Putin for 8 years.  Somehow this is Republican
slb42jcb|HuffPostBlog|0.4215|0.16|0.556|0.285|Why Hillary Lost: The Great American Lie https://t.co/mwvOaUzCDN via @HuffPostBlog
slb42jcb|huffingtonpost|0.4215|0.16|0.556|0.285|Why Hillary Lost: The Great American Lie https://t.co/mwvOaUzCDN via @HuffPostBlog
MJBodary|twitter|-0.8687|0.521|0.479|0.0|"You are disgusting human waste, JefferyGuterman.Hillary Clinton is a liar and a crook!#shameful https://t.co/g9zzvEYhMp"
LaborFAIL|GaetaSusan|-0.8594|0.399|0.498|0.103|"RT @GaetaSusan: Dems, McCain &amp; Graham STOP spreading FAKE NEWS! Every Country hacked Hillary's Private Server! Blame Russia?? What about bl"
JenniPxox|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
lorilpeabody|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
nytrbpolitics|nola|-0.7184|0.353|0.647|0.0|Hillary Clinton attacks 'fake news' in post-election appearance on Capitol Hill - https://t.co/w2DrHaeqHi https://t.co/K8C12gNu2L
TigernBham|peterjhasson|-0.4836|0.239|0.761|0.0|@peterjhasson @KerryPicket @DailyCaller How many million$ did Hillary keep after losing???
paulbenedict7|twitter|-0.7906|0.364|0.636|0.0|#Obamastan's FBI: no need to prosecute Hillary's uranium deal; Obamastan's CIA: Putin is a #Trump lobbyist. Worse t https://t.co/lai9DuXZLi
jerry_field|CobyRayan|0.807|0.0|0.673|0.327|"RT @CobyRayan: @CNN @GovChristie Made great history supporting @realDonaldTrump,he don't need job now!he's busy with crooked Hillary#lockhe"
NECEXAM|umpire43|-0.4215|0.113|0.887|0.0|RT @umpire43: Before the SC shut down MI Recount. several hundred thousand Hillary votes disqualified as poll book and vote boxes did not m
orangeteletubby|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
wvufanagent99|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
jihoonsthighs|maItinerecords|0.4019|0.0|0.838|0.162|RT @maItinerecords: hillary clinton flew all the way to hong kong to support twice https://t.co/Dsmufj6Xes
jihoonsthighs|twitter|0.4019|0.0|0.838|0.162|RT @maItinerecords: hillary clinton flew all the way to hong kong to support twice https://t.co/Dsmufj6Xes
720Sloan|HankDaTank25|0.5719|0.0|0.773|0.227|@HankDaTank25 @YouTube Hank i respect you but by that logic we should forgive Hillary for rigging the democrat primary
Kicker_Mom|TimOBrien|0.0|0.0|1.0|0.0|@TimOBrien @brianstelter Thought you were talking about Hillary for a moment
marlowstephens|twitter|-0.3612|0.116|0.884|0.0|"Hillary, Obama and SNL are clutching at straws. Their lazy assumptive attitude has bitten them on the rear end. https://t.co/Q2Xryo2Tcu"
CpturCre8Studio|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
HPLovecraft10|sbpdl|-0.5994|0.163|0.837|0.0|"RT @sbpdl: At this point, it's obvious the deep state is trying to instigate a civil war in USA over pro-Globalism Hillaryhttps://t.co/qOo"
sammy27932003|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
stuckin_mud|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
jwaters142|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
Patrioticgirl86|FreedomChild3|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
Patrioticgirl86|t|0.0|0.0|1.0|0.0|RT @FreedomChild3: HILLARY PLEADS TO DISMISS BENGHAZI LAWSUIThttps://t.co/5VxZ989pFd#BenghaziMatters #WakeUpAmerica https://t.co/uE4mKpX4
scott_stalker2|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
MoniqueCook20|umpire43|0.0|0.0|1.0|0.0|RT @umpire43: In Millwaukee day 5 of recount Hillary had 356000 votes thrown out for Fraud.Boxes in Millwaukee did not match poll books RUS
SireWilliamN|kashanacauley|-0.4767|0.205|0.795|0.0|RT @kashanacauley: It's a shame Hillary didn't connect with white Russian working class voters.
NPete2|Maldoduardo|0.0|0.0|1.0|0.0|RT @Maldoduardo: @DonaldsAngel @NPete2 @asamjulian @LindaSuhler @mitchellvii @Cernovich @JackPosobiec U suppose Hillary thinks it's #Fakene
1isten_up|PolitixGal|0.4404|0.0|0.756|0.244|RT @PolitixGal: Assessment of Hillary by her good friend... https://t.co/Wjdmabk7CF
1isten_up|twitter|0.4404|0.0|0.756|0.244|RT @PolitixGal: Assessment of Hillary by her good friend... https://t.co/Wjdmabk7CF
dcbdbc770706431|twitter|-0.6334|0.436|0.319|0.246|One more that's dumber is Hillary loser supporters crying like babies! https://t.co/9gC9Hmxugx
decook1961|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
DorAnnCecil|LindaSuhler|0.6523|0.0|0.835|0.165|RT @LindaSuhler: Only credible link to Russia is Hillary's -- who made herself RICH when she transferred 20% of our uranium to Putin...FOR
MiaEvan30311368|chuckie_chopper|0.0|0.0|1.0|0.0|RT @chuckie_chopper: @BreitbartNews @AJDelgado13 Hillary gave Russia US URANIUM and democrats claim Russia made @realDonaldTrump president?
Yougarte|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
Tamaraciocci|kylegriffin1|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
Tamaraciocci|theatlantic|-0.6597|0.293|0.707|0.0|RT @kylegriffin1: The Dangerous Myth That Hillary Clinton Ignored the Working Class @TheAtlantic https://t.co/bzCbt0iaXD https://t.co/Waam
frostdeeds|Online_Gangsta_|0.2023|0.136|0.679|0.185|@Online_Gangsta_ @justinhendrix @realDonaldTrump No it clever. Hillary's Goldman sachs connection is by money
bonniemurphy|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@AllenWest: ""It was President Obama, along with Hillary Clinton, that came up with the 'Russian reset button.'"" @JudgeJeanine"
Chlanandria|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
georgid63|bruce_arthur|0.7184|0.0|0.769|0.231|RT @bruce_arthur: Fun: imagine Hillary was elected with Russian help and gave donors cabinet posts and kept the Clinton Foundation and went
imnotheguy4you|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
USA4_Americans|usaforamericans|0.0|0.0|1.0|0.0|Trump: Bill Met AG Lynch on Jet to Offer Re-Appointment in a Hillary Clinton Admin https://t.co/LmSKiePOMb https://t.co/Dl5WvrXfV1
TrumpClaus|twitter|0.2732|0.145|0.617|0.238|Santa wishing #America a Merry Christmas &amp; #Hillary a long prison term at Trump Star Hollywood Ca. #MAGA https://t.co/pR32mmy9jB
Vote_American|Vote_American|-0.4926|0.285|0.715|0.0|@Vote_American Hillary should be Tried &amp; Convicted of Treason!
whatstherukkus|adamjohnsonNYC|0.4939|0.111|0.641|0.248|@adamjohnsonNYC Putin definitely gave Hillary the lowest favorable ratings of any candidate to ever run for the presidency.
MickeyJohnson07|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
keithingram214|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
_bigchee|ericgarland|0.6369|0.0|0.826|0.174|"RT @ericgarland: Hillary, for her part, gives a brief and all-too-calm speech and goes hiking. Probably the best move on the board."
drapes_vince|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
ladyleyn|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
t_ruggeri|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Tis4Ta|waitingroom8008|-0.4019|0.124|0.876|0.0|RT @waitingroom8008: things that are also true:1. Dems insisted that Hillary's FBI case wouldn't sway voters2. Hillary deserved to lose h
Proud1American|Stevenwhirsch99|-0.7088|0.257|0.743|0.0|@Stevenwhirsch99 @BooBreeze Using Clinton Foundation to hide foreign donations to Hillary's campaign was genius in a sinister kind of way!
NECEXAM|umpire43|0.0|0.0|1.0|0.0|RT @umpire43: In Millwaukee day 5 of recount Hillary had 356000 votes thrown out for Fraud.Boxes in Millwaukee did not match poll books RUS
_J32P_|HAWofPA|-0.8453|0.363|0.637|0.0|@HAWofPA Anyone paying attention hated Hillary LONG before a DNC insider leaked information. I notice Dems don't care about WaPo influence
Pooky_LoveRebel|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
alicewetterlund|matthewamiller|0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
alicewetterlund||0.0|0.0|1.0|0.0|RT @matthewamiller: It will be news to Hillary Clinton that the FBI will not draw inferences about things it can't prove in court. https://
mabian|HAGOODMANAUTHOR|-0.6808|0.219|0.781|0.0|RT @HAGOODMANAUTHOR: Hillary lost. Get over it establishment Democrats. You told Bernie voters to get over it. And you actually cheated Ber
jenmelton1976|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
jenmelton1976|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
ambitjournal|torontosun|-0.128|0.28|0.518|0.202|Hillary loved fake news  until she lost | Guest Column | World | News | Toronto https://t.co/z3T8xDO2YT
Txwench|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
RamBoPirate|xebec78|-0.5994|0.17|0.83|0.0|"RT @xebec78: @LeahR77 Hillary wanted to import 100k of them...must have been part of her master ""war on women"" plan..."
danmadio|nypost|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
danmadio|t|0.0772|0.111|0.766|0.123|RT @nypost: Hillary Clinton and her supporters spent twice as much as Donald Trump on her losing presidential campaign https://t.co/kPyf4Ns
Coach_For_LIfe|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
bbschumann|nia4_trump|-0.7096|0.258|0.742|0.0|RT @nia4_trump: Hillary blames Russia &amp; #FakeNews for her lossReality Check it was the Scandals Corruption Collusion &amp; Divisivenesshttps:
SnowMaylar|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
SnowMaylar|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
AriJameson|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
plz_think_1st|DaysOfTrump|-0.5994|0.196|0.804|0.0|"RT @DaysOfTrump: #AmericaFirst Patriots inside USgov are waging a civil war w international socialists (Hillary, Soros..) that have infiltr"
vipertoxin|youtube|0.2577|0.0|0.865|0.135|&gt;&gt; HILLARY WONT EVEN HAVE MAJORITY OF VOTES ONCE THE DUST CLEARS - YouTube https://t.co/qwS21s7WKT
ElaineCarlisl1|ElaineCarlisl1|0.7284|0.0|0.494|0.506|RT @ElaineCarlisl1: WIN BIG HILLARY!! https://t.co/2zXmCrSd2i
ElaineCarlisl1|twitter|0.7284|0.0|0.494|0.506|RT @ElaineCarlisl1: WIN BIG HILLARY!! https://t.co/2zXmCrSd2i
Richey4Fun|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
TroncaleJoseph|nia4_trump|0.0|0.0|1.0|0.0|RT @nia4_trump: Watch Hillary LIE during her SoS confirmation hearing. #ClintonCash #UraniumOne The RUSSIANS #ClintonFoundationhttps://t
Trillion3|CNNHeroes|0.0|0.0|1.0|0.0|@CNNHeroes @CNN https://t.co/kRF9EM73lH https://t.co/IHVrUxmhWm
Trillion3|thegatewaypundit|0.0|0.0|1.0|0.0|@CNNHeroes @CNN https://t.co/kRF9EM73lH https://t.co/IHVrUxmhWm
Scoote429143203|MissLizzyNJ|0.0|0.0|1.0|0.0|@MissLizzyNJ Oh Shush about Hillary! She has said nothing.
OTMOPTIONTWIT|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
OTMOPTIONTWIT|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
TheRavenxx|FratboyMarxist|0.3182|0.0|0.859|0.141|RT @FratboyMarxist: @fabucat @BlackAutonomist @angelsavant Hillary supported outright coups in countries overturning elected results (Hondu
atkinastarling|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
Vanila_Flav|GaetaSusan|-0.8594|0.399|0.498|0.103|"RT @GaetaSusan: Dems, McCain &amp; Graham STOP spreading FAKE NEWS! Every Country hacked Hillary's Private Server! Blame Russia?? What about bl"
VieuxBourru|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
EcuadorDeb|LPDLakeland|0.2023|0.137|0.637|0.225|"@LPDLakeland @Molon_Labe_Libs @1Kimsey @DineshDSouza Also, Obama can pardon Hillary, but there's no one to pardon Obama."
EmilyWA98498|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
scott_stalker2|asamjulian|-0.6159|0.285|0.611|0.104|RT @asamjulian: Funny watching libs cry about Russian interference (w/ no evidence) that didnt care at all about Hillarys MANY foreign i
CyndiLeeJ|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
CyndiLeeJ||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
Basilswiss|twitter|0.4404|0.0|0.734|0.266|"Thanks to Angela Merkel, Hillary Clinton, and Obama. https://t.co/JKVz1gF2bV"
jennifer4nm|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
KlinekeH50|LeahR77|0.0|0.0|1.0|0.0|"RT @LeahR77: Darn Those #RussianHackers If Only Libs Could Have Kept Hillary's Corruption, Fixing Primaries, &amp; Media Collusion Private She"
Rockprincess818|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
7brown30_06|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
TrinityNYC|t|0.0|0.0|1.0|0.0|https://t.co/FE3kumenP9CNN
UGA3949|FrankLuntz|-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
UGA3949||-0.1531|0.078|0.922|0.0|"RT @FrankLuntz: Did Russia also hack Hillary's campaign calendar and delete all her stops in rural Wisconsin, Penn., and Michigan?https:/"
conservogirl|asamjulian|0.7269|0.0|0.775|0.225|RT @asamjulian: How many months did the democrats have to investigate the source of Podestas email hacking? Funny they only care after Hil
altg03|twitter|0.7579|0.0|0.381|0.619|except she loves Hillary lol https://t.co/qD1o8PvHzw
statefarm2005|CNN|-0.705|0.328|0.672|0.0|"@CNN Hillary may have been reckless with her emails, but Trump is much worser."
Carlapaul18|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
kthedefused|MarkDice|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
kthedefused|youtube|-0.5411|0.179|0.821|0.0|RT @MarkDice: Hillary Clinton Wasted 1.2 Billion Dollars on Her Presidential Campaign!    Here's the Report:  https://t.co/8L8KaEbUzR http
WayneABryant|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
DragonTat2|KatieWagnerFox|0.3818|0.134|0.634|0.231|"RT @KatieWagnerFox: Seth Rich narc'd DNC emails because of cheating in Primary to promote Hillary. #SethRich, ultimate Bernie Bro, RIP. #"
jenmelton1976|MMsharbono|0.0|0.0|1.0|0.0|"RT @MMsharbono: Following their role model, Hillary. https://t.co/ShARZ1GtDw"
jenmelton1976|twitter|0.0|0.0|1.0|0.0|"RT @MMsharbono: Following their role model, Hillary. https://t.co/ShARZ1GtDw"
saveusrepublic2|WayneDupreeShow|-0.2023|0.217|0.664|0.119|"RT @WayneDupreeShow: There's no PROOF Russia hacked anything, let's be serious. The same media who said Hillary was winning in the polls is"
TonyWalker02|bfraser747|0.0129|0.19|0.617|0.193|"RT @bfraser747:  #ThanksObama You accomplished UR clear mission Stop blaming #RussianHackers &amp; #FoxNews#Hillary was a nightmare,  but"
strange_wulf132|LucidHuricane|0.7184|0.0|0.75|0.25|RT @LucidHuricane: The #UK has welcomed the trash of humanity into their country with open arms.  Hillary wanted this for USA. Thank god fo
JoanneFralin|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
Pas3652Paula|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
AmericanMom2|JudicialWatch|0.0|0.0|1.0|0.0|RT @JudicialWatch: In this country our leaders are bound by the rule of law. Hillary Clinton must be held accountable for her actions.http
MonlcaBabyyyy|ImBluetrek|-0.6402|0.246|0.754|0.0|RT @ImBluetrek: Donald Trump faked being upset with Hillary's emails. He does not care about Putin's Hackers https://t.co/9HwXKNP3Dx
MonlcaBabyyyy|twitter|-0.6402|0.246|0.754|0.0|RT @ImBluetrek: Donald Trump faked being upset with Hillary's emails. He does not care about Putin's Hackers https://t.co/9HwXKNP3Dx
sewingsandra|manny_ottawa|-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
sewingsandra||-0.3412|0.107|0.893|0.0|RT @manny_ottawa: How did even 1 person vote for Hillary.I can understand the deceased voting for her they didn't know better. https://t.c
PensiveTM|mtracey|-0.7728|0.317|0.605|0.078|"RT @mtracey: @bhking03897 @kthalps The problem lies in Hillary setting up a private server, lying about it, and running despite severe lega"
wyodebbie|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: People weren't concerned about Russia when Hillary was selling them US uranium.#MAGA
Eliz_Hightower|cjsienna55|-0.5267|0.159|0.841|0.0|RT @cjsienna55: @TheLiePolitic @TheDonaldNews  I tell you people on the inside had to be disgusted with what Hillary was doing.
HeddRoxx|usacsmret|0.1232|0.0|0.928|0.072|"RT @usacsmret: ""FakeNews"" doesn't explain Hillary's loss, but it does describe the media's coverage of Obama these past eight years."
Anzers|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
steveinashland|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
MiaEvan30311368|JodyCoyote12|-0.6908|0.231|0.769|0.0|"RT @JodyCoyote12: @NJTrumpWarrior @BreitbartNews No, it's a last ditch attempt by elites to get Hillary's corrupt ass into the WH where she"
TheOnly313Girl|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
kenwheaton|notjessewalker|0.0|0.0|1.0|0.0|"RT @notjessewalker: Evergreen line: ""The Obama administrationperhaps anticipating a Hillary Clinton presidencysupported these changes"" ht"
KarenSeasly|umpire43|0.5107|0.101|0.645|0.253|"RT @umpire43: BOMBSHELL VIDEO : The NSA, not Russia, HACKED the DNC to Help Derail a Hillary Presidency https://t.co/RLMA0vm53R"
KarenSeasly|linkis|0.5107|0.101|0.645|0.253|"RT @umpire43: BOMBSHELL VIDEO : The NSA, not Russia, HACKED the DNC to Help Derail a Hillary Presidency https://t.co/RLMA0vm53R"
Lori_Bardsley|RichardGrenell|0.4019|0.11|0.705|0.185|RT @RichardGrenell: I'd love to know how the Russians got Hillary to ignore union workers in the Midwest.
AU_bebe|TrumpCard555|0.8134|0.114|0.492|0.394|RT @TrumpCard555: Agree @Rosechristenbe1 they were so confident #hillary would win &amp; panicked since. Hundreds-thousands #Illegals brought h
Truest_Thoo|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
SeesEarth|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
SeesEarth||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
TRUMPIS4US|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
scott_stalker2|MStuart1970|0.4199|0.0|0.866|0.134|RT @MStuart1970: RUSH: While Trump Tours To Thank America... Look What The Hildebeast Is Up To! https://t.co/iPK5Cxrk7M via @Doug_Giles#T
scott_stalker2|clashdaily|0.4199|0.0|0.866|0.134|RT @MStuart1970: RUSH: While Trump Tours To Thank America... Look What The Hildebeast Is Up To! https://t.co/iPK5Cxrk7M via @Doug_Giles#T
rmack2x|halsteadg048|0.0|0.0|1.0|0.0|RT @halsteadg048: Hillary Clinton Takeover of the USA https://t.co/WyvI6OVBrT PROOF By Dr Pieczenik Counter-Coup Who Worked w/ Julian To St
rmack2x|youtube|0.0|0.0|1.0|0.0|RT @halsteadg048: Hillary Clinton Takeover of the USA https://t.co/WyvI6OVBrT PROOF By Dr Pieczenik Counter-Coup Who Worked w/ Julian To St
shrewst|KatieWagnerFox|0.3818|0.134|0.634|0.231|"RT @KatieWagnerFox: Seth Rich narc'd DNC emails because of cheating in Primary to promote Hillary. #SethRich, ultimate Bernie Bro, RIP. #"
Trinidadiyon|France4Hillary|0.34|0.082|0.786|0.132|"RT @France4Hillary: #Hillary lost 4 states (FL, MI, WI, PA) by ~1 point. If not for Russia/Comey, she'd have won them all. WE NEED A #REVOT"
Lena_D_Sarcast|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
Alllwftopic|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
kelly77_ryan|LadyPatriot2000|-0.4939|0.158|0.842|0.0|RT @LadyPatriot2000: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #tcot https://t.co/1wlS
kelly77_ryan|t|-0.4939|0.158|0.842|0.0|RT @LadyPatriot2000: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #tcot https://t.co/1wlS
Raelyk|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
Steven_Strauss|DustinGiebel|-0.4019|0.172|0.828|0.0|RT @DustinGiebel: Hillary hacked the DNC because Trump was hogging all the attention.  #BoltonFalseFlagExcuses
TheOxyCon|NotJoshEarnest|0.0|0.0|1.0|0.0|RT @NotJoshEarnest: Hillary tried to go to Wisconsin and Michigan but the Russians kept hacking her plane back to California and New York
DrJillJoyce|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
DrJillJoyce||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
EightyNine10|eightynine10studios|0.5319|0.0|0.791|0.209|HILLARY CLINTON IS THROWING A PARTY -- YOU WON'T BELIEVE THE REASON WHY - https://t.co/PGb9pDUqOR https://t.co/DI2QSgU2qW
pyowac1|thehill|-0.7579|0.306|0.694|0.0|@thehill Only the gullible believe that Hillary is guilty of all that she is accused of. Most of it unfounded
CpturCre8Studio|StevePieczenik|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
CpturCre8Studio|t|-0.608|0.296|0.529|0.175|RT @StevePieczenik: luv #podestaspizza reference HELL o #America knows the scoop #Hillary have some dignity LEAVE #pizzagate https://t.co/w
JamesRitch1|Duane106|-0.7003|0.266|0.734|0.0|"RT @Duane106: After She Criticized Hillary, 'Morning Joe' Anchor Says NBC Got a Disturbing Call from Clinton Campaign... https://t.co/q6TiV"
JamesRitch1|t|-0.7003|0.266|0.734|0.0|"RT @Duane106: After She Criticized Hillary, 'Morning Joe' Anchor Says NBC Got a Disturbing Call from Clinton Campaign... https://t.co/q6TiV"
username__111|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: I repeat: I laid out what was going on with Russian campaign, based on leaks from European intel, before election: http"
dreamerbeast|FrankConniff|-0.9136|0.394|0.606|0.0|"RT @FrankConniff: Don't give me that ""Hillary was a bad candidate"" bullshit. Real-life Bond villains plotted against her and she still got"
Denicebrown2000|KailiJoy|0.0|0.0|1.0|0.0|"RT @KailiJoy: Anyway. You can expect that I'll be talking about Hillary Clinton, the president who should have been, for the next four year"
gerfingerpoken2|americanthinker|-0.5106|0.202|0.798|0.0|#Benghazi Mom Patricia Smith Targets Serial Liar Hillary https://t.co/KVO6ImiEzS - American Thinker - #PJNET 999 - https://t.co/Jiwbz2JGaU
annie5133|DustinGiebel|-0.4019|0.172|0.828|0.0|RT @DustinGiebel: Hillary hacked the DNC because Trump was hogging all the attention.  #BoltonFalseFlagExcuses
WVaChris2|dcexaminer|0.7707|0.0|0.767|0.233|@dcexaminer Is this the same Silver who said Hillary was a sure bet to win on Election Day despite know if FBI investigation? Sour Grapes!!
musthavebeenme|PhilipRWFG|0.3527|0.109|0.724|0.167|RT @PhilipRWFG: @politico So he's saying Obama hacked Hillary and pretended to be Russia so that Trump could win? Huh?
Mster_Carpentr|LibertyLivesHer|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
Mster_Carpentr|vivaliberty|-0.3818|0.206|0.794|0.0|RT @LibertyLivesHer: Hillarys Losing Campaign Cost a Record $1.2 Billion - #ClintonCash https://t.co/hNgphruaE7
karenmi49109968|peterjhasson|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
karenmi49109968|dailycaller|-0.4939|0.158|0.842|0.0|RT @peterjhasson: Hillary Donors Could Have Fed 6 Million Hungry Children For A Year With Wasted Campaign Money https://t.co/a9yjWWX9eF via
casualhypocrite|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
catwahler|gerfingerpoken2|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
catwahler|floppingaces|0.0|0.0|1.0|0.0|"RT @gerfingerpoken2: Trump Defends Life, Hillary Defends Partial Birth Abortion - Flopping Aces - https://t.co/3vfWU1mTTb #MAGA #PJNET http"
MoniqueCook20|TweetingYarnie|-0.4599|0.228|0.616|0.156|RT @TweetingYarnie: I never get tired of reading how arrogant and wrong Hillary Clinton's campaign was despite warnings that she could loos
ghostofanation|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
ghostofanation|t|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
azjennytobin|redsteeze|0.0|0.0|1.0|0.0|RT @redsteeze: Russia wanted Trump. You know who else wanted Trump? Hillary &amp; our media. All three got what they wanted.
npnikk|npnikk|-0.1396|0.137|0.75|0.113|"RT @npnikk: Joe Scarborough It wasnt fake news."" Hillary Clinton Cost Hillary Clinton the Election, Not Fake News. https://t.co/fzcvbyI"
npnikk|t|-0.1396|0.137|0.75|0.113|"RT @npnikk: Joe Scarborough It wasnt fake news."" Hillary Clinton Cost Hillary Clinton the Election, Not Fake News. https://t.co/fzcvbyI"
PRrodLA|stacyherbert|-0.3182|0.108|0.892|0.0|RT @stacyherbert: Pew says Hillary lost big with middle class voters | I say: exactly income brackets paying full Obamacare premiums https:
kelly77_ryan|IdiotDems|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
kelly77_ryan|t|-0.4939|0.158|0.842|0.0|RT @IdiotDems: Hillary Donors Could Have Fed 6 Million Hungry Children For a Year With Wasted Campaign Cash - #CrookedHillary https://t.co/
mattlast84|StefanMolyneux|-0.4588|0.125|0.875|0.0|RT @StefanMolyneux: Cant wait for Dem investigation to figure out how Russian hackerz (TM) forced Hillary to take millions in Saudi money.
ElDon78|twitter|-0.5255|0.298|0.702|0.0|What&gt; Bolton is wrong. Hillary did the hacking! https://t.co/Out6NltZJc
queenofsoul62|KellyannePolls|-0.783|0.261|0.652|0.087|"@KellyannePolls why you guys still at Hillary, election over we doomed to hell judge not lest he be judged he without sin cast first stone."
TommyVape|LindaSuhler|0.4404|0.0|0.847|0.153|RT @LindaSuhler: A good time to mention Hillary Clinton's REAL link to Russia...#RussianHackingShe transferred our uranium to Putin...FOR
lkdavolos|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
lkdavolos|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
danfelix82|HeideggerFan|0.4588|0.0|0.842|0.158|@HeideggerFan @Lglwry @justinhendrix @realDonaldTrump @PolitiFact yet crickets from you on the liberal media reporting to benefit Hillary...
wclay1|ScottyLiterati|-0.296|0.091|0.909|0.0|RT @ScottyLiterati: Hillary dropped this exact same info about Russia in front of 66 million viewers in October. But I guess no one listene
GretchenInOK|asamjulian|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
GretchenInOK|realclearpolitics|-0.3612|0.152|0.848|0.0|RT @asamjulian: Priebus: The Russians Didn't Force Hillary Clinton To Ignore Wisconsin and Michigan  https://t.co/IFOVeb3LXd
Kimberley1222|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
bbeennny|peddoc63|0.1531|0.084|0.812|0.104|RT @peddoc63: Do you care that Hillary sold 20% of our Uranium to Russians? Or that Obama lied to pass Iran Deal &amp; Obamacare &amp;that he paid
rodsandguitars|politico|-0.6966|0.229|0.771|0.0|@politico Remember IRS targeting? Remember DOJ Contempt of Congress? Remember Benghazi coverup? Remember Hillary's Nuclear Material Deal?
erincowgill|Craigipedia|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
erincowgill|twitter|-0.6369|0.208|0.792|0.0|"RT @Craigipedia: Remember all the geniuses who voted against Hillary because they hated ""the Clinton Dynasty""? https://t.co/rwJ4K9dlmO"
MargaretMcgui16|Ian56789|-0.4588|0.13|0.87|0.0|RT @Ian56789: Remember when Russian Hackers forced Hillary to wipe her server after being served with a Congressional Sub Poena to preserve
rebelgirl1776|RepStevenSmith|0.0772|0.0|0.939|0.061|RT @RepStevenSmith: Want to hear about what Hillary did in Libya from a real journalist? @wikileaks Julian Assange explains it in 2 minutes
kimberlymontse1|twitter|0.8689|0.0|0.597|0.403|They increase #ProfitCare business though.. thanks to Hillary &amp; friends like #FDA #CDC working to COVER UP the fact https://t.co/56hk8obyRP
TruthqueenVA|Change|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/RZBqJtPhx0 via @Change
TruthqueenVA|change|-0.296|0.196|0.804|0.0|You Can Stop Trump on December 19 https://t.co/RZBqJtPhx0 via @Change
NPete2|DaysOfTrump|-0.5994|0.196|0.804|0.0|"RT @DaysOfTrump: #AmericaFirst Patriots inside USgov are waging a civil war w international socialists (Hillary, Soros..) that have infiltr"
TheBeijingKing_|jasonroeder|-0.4215|0.149|0.851|0.0|"RT @jasonroeder: Too late to point fingers, but did Hillary make even ONE campaign stop in Moscow?"
osoloco11|CronkiteSays|-0.3818|0.205|0.697|0.098|RT @CronkiteSays: REAL NEWSWe've completed an extensive analysis into why Hillary lost and have determined Hillary caused Hillary to lose
RealNaylorSmall|TrumpSuperPAC|-0.7772|0.244|0.756|0.0|RT @TrumpSuperPAC: We came close to the apocalypse with this raving lunatic! #Hillary wants to censor all media! Who's the Nazi now? https:
CROWENATION2016|TweetingYarnie|-0.4599|0.228|0.616|0.156|RT @TweetingYarnie: I never get tired of reading how arrogant and wrong Hillary Clinton's campaign was despite warnings that she could loos
TypicalHenshiri|LibyaTopTweets|0.0|0.0|1.0|0.0|RT @LibyaTopTweets:                     htt
saket016|MissLizzyNJ|0.2732|0.0|0.896|0.104|"RT @MissLizzyNJ: Hillary Clinton, who accepted millions from Saudi Arabia &amp; Qatar, is suddenly concerned about foreign governments influenc"
constantino_sam|pinterest|0.1598|0.171|0.565|0.263|HILLARY FOR PRESIDENT? You F**CKING  Kidding Me? ANTI HILLARY Funny Bumper Stick https://t.co/VkKQtKj3gV
patlinetweet|FoxNews|-0.6901|0.222|0.778|0.0|"RT @FoxNews: .@GovMikeHuckabee: ""It wasn't the Russians that beat them. It was a lack of ideas. It was Hillary being a very poor candidate."
katherinejnowak|teeg_dougland|0.3491|0.053|0.842|0.106|@teeg_dougland @neeratanden 50. making hillary dab on ellen &amp; appear on broad city but not apologize for hurting black comm in 08 &amp; 1st lady
meezer16|DaysOfTrump|-0.5994|0.196|0.804|0.0|"RT @DaysOfTrump: #AmericaFirst Patriots inside USgov are waging a civil war w international socialists (Hillary, Soros..) that have infiltr"
maattlyons|WalshFreedom|0.5859|0.0|0.84|0.16|"RT @WalshFreedom: If there was evidence that the Russians helped Hillary win, my fellow conservatives would be yelling for an investigation"
Alllwftopic|ericgarland|0.8761|0.0|0.654|0.346|"RT @ericgarland: I'm from Vermont and have known Bernie forever, so I'm very surprised, but everyone kinda likes it. Hillary wins anyhow."
khelfrich08|LisaToddSutton|0.6114|0.0|0.688|0.312|"@LisaToddSutton @KellyannePolls lol, okay. Hillary is the president-elect! Time to take your medication."
Williamwvaughn|bessbell|-0.5574|0.217|0.709|0.075|@bessbell @realDonaldTrump joking right? He was elected because Hillary and the liberals have no message and failed polices. Give me a break
Phyllis28333|Lrihendry|-0.5848|0.147|0.853|0.0|"RT @Lrihendry: If Russia is the enemy, why didn't anyone look into why Hillary sold 20% of our uranium to them! #FakeNewsChallenge @realDon"
Shishu40011004|Sterlingartz|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
Shishu40011004|motherjones|0.4215|0.0|0.865|0.135|RT @Sterlingartz: hillary clinton's lead in the popular vote swells to nearly 2.7 million and 48% ... https://t.co/ro7TGgtxEW https://t.co/
_bigchee|ericgarland|-0.0516|0.101|0.806|0.093|"RT @ericgarland: And now, the target for electoral mischief is enormous. Hillary is the most known quantity in America, with huge backstory."
dakotahsmom6|datrumpnation1|0.0|0.0|1.0|0.0|RT @datrumpnation1: Look who is behind the Russian CIA story:1. Washington Post2. Obama3. Schumer 4. McCain &amp; Lindsay Graham5. Hillary
ErickaJacobs123|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
