User|Original_User/Web|Compound|Negative|Neutral|Positive|Tweet
mapocoloco|nytimes|0.4767|0.0|0.853|0.147|"RT @nytimes: Donald Trump indicated that, as president, he would take the daily intelligence briefing ""when I need it"" https://t.co/3V8bqwm"
mapocoloco|t|0.4767|0.0|0.853|0.147|"RT @nytimes: Donald Trump indicated that, as president, he would take the daily intelligence briefing ""when I need it"" https://t.co/3V8bqwm"
DonMcKenzie|Delo_Taylor|-0.4404|0.14|0.86|0.0|RT @Delo_Taylor: I was never 100% on board with Bernie &amp; some of his Stans may have been obnoxious but they did have a plan for stopping Tr
rappahannockmag|JohnWDean|-0.6597|0.188|0.76|0.052|"RT @JohnWDean: Notwithstanding Trump's efforts to kill this, there are a few real Americans in the US Senate who want answers: https://t.co"
rappahannockmag|t|-0.6597|0.188|0.76|0.052|"RT @JohnWDean: Notwithstanding Trump's efforts to kill this, there are a few real Americans in the US Senate who want answers: https://t.co"
schober_lisa|arnonmishkin|-0.3818|0.133|0.867|0.0|@arnonmishkin @Martina @Bencjacobs Trumps father had Alzheimer's.  Trump is showing signs himself.  He is being manipulated by Russia.
serge_poznanski|ft|0.34|0.0|0.876|0.124|"FT: Trump puts four-decade old ""One China"" policy in play: Trumps position is you can trade anything  https://t.co/sqhZdwbYkr"
thalsey51|DCClothesline|-0.4588|0.232|0.67|0.098|Secret CIA Assessment Story About Russia Helping Trump is Fake News Youve Been Warned About https://t.co/uMG6yQmixc via @DCClothesline
thalsey51|linkis|-0.4588|0.232|0.67|0.098|Secret CIA Assessment Story About Russia Helping Trump is Fake News Youve Been Warned About https://t.co/uMG6yQmixc via @DCClothesline
sweettea4me925|amjoyshow|0.0|0.0|1.0|0.0|RT @amjoyshow: Trump advisers with Russian ties https://t.co/hISlPTqQ2m via @amjoyshow
sweettea4me925|msnbc|0.0|0.0|1.0|0.0|RT @amjoyshow: Trump advisers with Russian ties https://t.co/hISlPTqQ2m via @amjoyshow
lord_rosenberg|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
semirabella|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
semirabella||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
puppy_training_|twitter|0.0|0.0|1.0|0.0|#WolrdNewsNew York TimesTrump Suggests Using Bedrock China Policy as Bargaining ChipNew York TimesPresident-ele https://t.co/dMTHtcInKe
LetsSeeLife|ObamaMalik|0.4019|0.0|0.828|0.172|RT @ObamaMalik: Let us support those who were in the fox hole with Mr.Trump.
TerrySoileau|ABCPolitics|-0.4215|0.192|0.808|0.0|"RT @ABCPolitics: Poll shows public skeptical over key Trump proposals, from cutting environmental regulations to repealing Obamacare https:"
LSoudek|CaptainsLog2016|0.1531|0.097|0.784|0.119|RT @CaptainsLog2016: Donald Trump is pretty upset because Navy didn't winHe was going to root for ArmyBut then he found out they were n
WLSTONE1|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
WLSTONE1||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
AppleCupBlues|twitter|0.8402|0.0|0.64|0.36|"""...the combined wealth of Trump's prospective cabinet tops $14 billion  more than 30 times greater than that of e https://t.co/jnpVl5HOmi"
OliviaAllenC|breitbart|-0.4767|0.181|0.819|0.0|"Rand Paul: Unrealistic, Unfair to Expect Trump to Sell All of His Businesses https://t.co/Epq0lgPFK8 https://t.co/B530oW4tyM"
intl_traveller|davidfrum|0.7351|0.0|0.754|0.246|"RT @davidfrum: US intelligence community: Russia acted to install Trump. 18 months from now, there wont be a US intelligence community wor"
AnonBruja|McClatchyDC|0.5859|0.0|0.826|0.174|"RT @McClatchyDC: Since his election win, Trump has talked to Putin more than any other world leader https://t.co/mLBJ0589N3 https://t.co/QN"
AnonBruja|mcclatchydc|0.5859|0.0|0.826|0.174|"RT @McClatchyDC: Since his election win, Trump has talked to Putin more than any other world leader https://t.co/mLBJ0589N3 https://t.co/QN"
eloinformada|franchosa|0.0|0.0|1.0|0.0|RT @franchosa: Empiezo a entender por qu gan Trump https://t.co/OhmRp3ubzc
eloinformada|twitter|0.0|0.0|1.0|0.0|RT @franchosa: Empiezo a entender por qu gan Trump https://t.co/OhmRp3ubzc
FactorsTalcott|yojudenz|0.6808|0.0|0.752|0.248|RT @yojudenz: Trump Is Planning on Giving Up a Presidential Luxury to Save 'Out of Control' Cost to Taxpayers https://t.co/HDaiBi20jR
FactorsTalcott|ijr|0.6808|0.0|0.752|0.248|RT @yojudenz: Trump Is Planning on Giving Up a Presidential Luxury to Save 'Out of Control' Cost to Taxpayers https://t.co/HDaiBi20jR
KarmaKittySays|V_of_Europe|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
KarmaKittySays|thegatewaypundit|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
OldBarbedWire|twitter|0.0|0.0|1.0|0.0|We hang on your every tweet Mr. Trump. https://t.co/GBkGFsCEco
gisellegrenier|cjcmichel|0.0|0.0|1.0|0.0|"RT @cjcmichel: Wife of Richard Spencer, alt-right figurehead, has translated writings of Alexander Dugin: https://t.co/x9jh55bO2V"
gisellegrenier|motherjones|0.0|0.0|1.0|0.0|"RT @cjcmichel: Wife of Richard Spencer, alt-right figurehead, has translated writings of Alexander Dugin: https://t.co/x9jh55bO2V"
EVIL_DAESH|dailystar|-0.8625|0.389|0.521|0.09|#US #China war is coming: World War 3 threat as China promises more nukes to 'prepare' https://t.co/ed43wPZcrR #WorldWar3 #NuclearWar #USA
KRCSmith62|MrDane1982|-0.25|0.14|0.755|0.104|RT @MrDane1982: At this point you look un-American while supporting Russia war with America. Donald Trump works for Putin not with him. htt
BourneInTexas|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
AlwaysAgnew|abbydphillip|-0.3724|0.118|0.882|0.0|"RT @abbydphillip: Trump on Fox News Sunday says he doesn't need daily intelligence briefings as POTUS because he's ""smart"" https://t.co/OUi"
AlwaysAgnew|t|-0.3724|0.118|0.882|0.0|"RT @abbydphillip: Trump on Fox News Sunday says he doesn't need daily intelligence briefings as POTUS because he's ""smart"" https://t.co/OUi"
RickySi16087724|shannonsbeau|0.6369|0.0|0.785|0.215|@shannonsbeau  I sure hope Trump watches His back side He's uncovering corruption that we would never of known if not for Him
baumsche|msn|-0.743|0.412|0.588|0.0|"Before Trump, there was a Muslim registry. It caught no terrorists https://t.co/QXHn9of1Gy"
Sciencereport36|itechpost|0.0772|0.0|0.894|0.106|What Future Awaits The Science Department Under Trump Administration? - iTech Post https://t.co/d5nbMFZTmx
B_Zamacona|reforma|-0.34|0.13|0.87|0.0|La comunidad de inteligencia de EU se alarm ante los comentarios y el rechazo de Donald Trump https://t.co/P7BzK25ytM
Zelidasquare|vermaak_martin|-0.6454|0.193|0.807|0.0|RT @vermaak_martin: @mitchellvii They have to stay the course as they have no choice If Trump did not win The media would start operating
rprez2012|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
NickRiccardi|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
NickRiccardi||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
MoMeldrum|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
zwwwara|amjoyshow|-0.4404|0.132|0.868|0.0|"RT @amjoyshow: Scott Dworkin (@FUNDER) started #TrumpLeaks documenting hundreds of Trump's Russian ties, which the #FBI has denied or not r"
mile_high_33|AndNowIWrite|0.3834|0.057|0.828|0.115|@AndNowIWrite how would you know when it's been your type in charge for last 8 yrs. trump will save this country and u idiots won't admit it
matometrump|trump|0.0|0.0|1.0|0.0|   livedoor https://t.co/qbstkpUtD1
Mr_Zues_1|DavidCornDC|0.6705|0.0|0.732|0.268|"@DavidCornDC A thought: Alec Baldwin,as trump,does intelligence briefings on SNL.trump will think he's giving the briefings to himself."
donkosin|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: When Obama used Dijon mustard, Fox attackd him 4 not using yellow mustrd (true) Yet they shrug when Trump says doesnt n"
Kirstycat1209|GusSent|0.6908|0.0|0.801|0.199|"RT @GusSent: Now calculate the value of all the free, excessive airtime for Trump by tv media--and realize the money was spent, just not by"
GalinaGalanos|bennydiego|0.0772|0.13|0.725|0.145|"RT @bennydiego: ""Nobody really knows"" except the entire scientific community. His ignorance is astounding. #climatechange https://t.co/f2yp"
GalinaGalanos|t|0.0772|0.13|0.725|0.145|"RT @bennydiego: ""Nobody really knows"" except the entire scientific community. His ignorance is astounding. #climatechange https://t.co/f2yp"
LKuehn4|kurteichenwald|0.5574|0.0|0.847|0.153|"RT @kurteichenwald: If Trump started getting praise 4  appointments from ISIS, do you think Fox News would start running stories about how"
KohenBrady|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
FilistineNow|nytimes|0.0|0.0|1.0|0.0|"#MedioOriente Boeing Seeks to Sell Planes to Iran, and the Deal to Trump https://t.co/2zRKNnIW6c #NYTIMES"
bluedevildavey|IslamismMap|-0.4215|0.177|0.823|0.0|"RT @IslamismMap: #MuslimBrotherhood's CAIR (https://t.co/TEMgYRfHfu) fears @GenFlynn, bc he believes #Islamism is existential threathttps:"
bluedevildavey|islamism-map|-0.4215|0.177|0.823|0.0|"RT @IslamismMap: #MuslimBrotherhood's CAIR (https://t.co/TEMgYRfHfu) fears @GenFlynn, bc he believes #Islamism is existential threathttps:"
CoryKCrabtree|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
CoryKCrabtree|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
partynauseous27|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
NewsLycaness19|frankrichny|-0.1603|0.064|0.936|0.0|"RT @frankrichny: By holding back RNC emails, Putin didn't just help install Trump in White House but has means to blackmail GOP to do his b"
Old96er1|keithlaw|0.0|0.0|1.0|0.0|@keithlaw @jnpaquet I heard that Trump really does poop his pants though.
goffmania|Noahpinion|-0.6124|0.263|0.647|0.091|"RT @Noahpinion: Prediction: Trump will push hard to kill alternative energy technology. After all, Russia is a petrostate... https://t.co/f"
goffmania|twitter|-0.6124|0.263|0.647|0.091|"RT @Noahpinion: Prediction: Trump will push hard to kill alternative energy technology. After all, Russia is a petrostate... https://t.co/f"
a_hundred_tacks|mattyglesias|0.4019|0.109|0.628|0.264|RT @mattyglesias: Trump pretending to dislike the network that hired a special stable of relentlessly pro-Trump pundits is egregious https:
Fernasteady|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
hwhlj321|BrettArends|0.5411|0.0|0.851|0.149|"RT @BrettArends: Hey, Netanyahu! If #Trump is such a friend of Jews, why does he hang out with Ann ""f---ing Jews"" Coulter?"
KimShirley123|pharris830|0.0|0.0|1.0|0.0|RT @pharris830: President Obama showing Trump around the Oval Office! https://t.co/pm8lVyGsFY
KimShirley123|twitter|0.0|0.0|1.0|0.0|RT @pharris830: President Obama showing Trump around the Oval Office! https://t.co/pm8lVyGsFY
StephanieMilli3|PrisonPlanet|-0.5574|0.261|0.739|0.0|RT @PrisonPlanet: Michael Moore: Something Crazy Could Happen to Stop Trump Becoming President - https://t.co/voVcYwLTJx https://t.co/WD0
StephanieMilli3|infowars|-0.5574|0.261|0.739|0.0|RT @PrisonPlanet: Michael Moore: Something Crazy Could Happen to Stop Trump Becoming President - https://t.co/voVcYwLTJx https://t.co/WD0
joh53293471|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
LE_Durfey|FT|0.34|0.0|0.882|0.118|"RT @FT: Trump puts four-decade old ""One China"" policy in play: Trumps position is you can trade anything  https://t.co/QEyRMK01nQ"
LE_Durfey|ft|0.34|0.0|0.882|0.118|"RT @FT: Trump puts four-decade old ""One China"" policy in play: Trumps position is you can trade anything  https://t.co/QEyRMK01nQ"
JLovrensky|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
Sciencesharenew|itechpost|0.0772|0.0|0.894|0.106|What Future Awaits The Science Department Under Trump Administration? - iTech Post https://t.co/VprQLvedXB
Patrioticgirl86|JrcheneyJohn|0.0|0.0|1.0|0.0|RT @JrcheneyJohn: The #FakeNews Media has been Neutered by Trump and they have become Irrelevant #TrumpEffect  https://t.co/8ArN8MrraK
Patrioticgirl86|twitter|0.0|0.0|1.0|0.0|RT @JrcheneyJohn: The #FakeNews Media has been Neutered by Trump and they have become Irrelevant #TrumpEffect  https://t.co/8ArN8MrraK
caitlinsloanx|charlymim|0.0|0.167|0.667|0.167|RT @charlymim: Why does my dad look like Donald Trump :-(  https://t.co/qRToKfj8q1
caitlinsloanx|twitter|0.0|0.167|0.667|0.167|RT @charlymim: Why does my dad look like Donald Trump :-(  https://t.co/qRToKfj8q1
KristaKaroFL|realDonaldTrump|0.3612|0.0|0.902|0.098|".@realDonaldTrump Trying to get Trump to read intel reports instead of watch tv, is like telling ur kids to do their homework on a weekend."
grandpooba5440|ActionTime|0.6739|0.0|0.799|0.201|RT @ActionTime: CIA: Russia Stole Presidency via Trump.US Electoral College Can WIN It Back #NotMyPresident #Resistance #Resist #RT https:/
grandpooba5440||0.6739|0.0|0.799|0.201|RT @ActionTime: CIA: Russia Stole Presidency via Trump.US Electoral College Can WIN It Back #NotMyPresident #Resistance #Resist #RT https:/
agrippa550|LindaSuhler|-0.5423|0.22|0.78|0.0|RT @LindaSuhler: The Silent Majority STOOD with Donald J. Trump and we shocked the world.Never underestimate pissed-off Patriots.#Presid
evelinekipping|HuffingtonPost|0.0|0.0|1.0|0.0|"RT @HuffingtonPost: Trevor Noah still can't figure out why Donald Trump calls China ""Jina"" https://t.co/qV216LQLMv https://t.co/lI5LkfdFpu"
evelinekipping|m|0.0|0.0|1.0|0.0|"RT @HuffingtonPost: Trevor Noah still can't figure out why Donald Trump calls China ""Jina"" https://t.co/qV216LQLMv https://t.co/lI5LkfdFpu"
KroekerTony|tazie34|0.4466|0.0|0.827|0.173|RT @tazie34: Traitors John McCain and Lindsey Graham JOIN DEMOCRATS to DELEGITIMIZE President-Elect Trump https://t.co/a0SzOaW8mx
KroekerTony|truthfeed|0.4466|0.0|0.827|0.173|RT @tazie34: Traitors John McCain and Lindsey Graham JOIN DEMOCRATS to DELEGITIMIZE President-Elect Trump https://t.co/a0SzOaW8mx
ShawnMorse_|GrrrGraphics|0.0|0.0|1.0|0.0|RT @GrrrGraphics: New #BenGarrison #Cartoon #NewBroom #Trump #Maga Sweep away the dirt/ #FakeNews ! more cartoons at https://t.co/Oj98iIxEA
ShawnMorse_|t|0.0|0.0|1.0|0.0|RT @GrrrGraphics: New #BenGarrison #Cartoon #NewBroom #Trump #Maga Sweep away the dirt/ #FakeNews ! more cartoons at https://t.co/Oj98iIxEA
JkFlower60|seankent|0.9179|0.0|0.536|0.464|"RT @seankent: Trump voters, does this seem like a legit reason for skipping intelligence briefings? Does it inspire confidence?   https://t"
JkFlower60||0.9179|0.0|0.536|0.464|"RT @seankent: Trump voters, does this seem like a legit reason for skipping intelligence briefings? Does it inspire confidence?   https://t"
oxfordtarheel|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: We CANT be split lib/conserv or GOP/Dem over Russia hack issue. This is an American issue. Trump can prove he is indepe
FMAlchemist|BillMoyersHQ|-0.6808|0.239|0.761|0.0|RT @BillMoyersHQ: To #Trump from Bill Moyers &amp; @MichaelWinship: No bribes in the form of tax cuts for big business. No backdoor deals. http
Figment_Imagine|twitter|0.0|0.0|1.0|0.0|But he's a white male who fawns over tRump. https://t.co/j9aXeayRhT
martycoultas|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
Libertarian896|slone|-0.5267|0.127|0.833|0.04|"RT @slone: YOU McCain are a ""matter of concern"" to Trump voters. YOU are a globalist pig who has helped destroy the US and the world. ENOUG"
Espormibien|bessbell|0.0|0.0|1.0|0.0|@bessbell @realDonaldTrump real Americans voted Trump!!  Not #clintonstench
pianodiva11|ClimateCentral|0.0|0.0|1.0|0.0|"RT @ClimateCentral: Trump's pick to run the Interior Department, Cathy McMorris Rodgers, has an extreme anti-environment voting record ht"
oufenix|TheGnudz|0.0516|0.089|0.813|0.098|RT @TheGnudz: @RachieBabe079 Why do you people keep giving Trump a pass when he's actually doing the very things you falsely accused Clinto
JenRothe|kurteichenwald|0.7089|0.0|0.772|0.228|"RT @kurteichenwald: Trump says: So smart doesnt need daily intel briefings, knows more about ISIS than military, knows tax code better than"
razzleberry_e|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
razzleberry_e|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
XMerc45|blaubok|0.47|0.096|0.652|0.252|RT @blaubok: When her election was 98% certain - Hillary assured Trump - the election isn't riggedWhen she lost - the election was rigged
TruthTeamOne|MrJamesonNeat|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
TruthTeamOne|t|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
georgebrown06|TheDailyEdge|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
georgebrown06|twitter|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
Aviationshare|usatoday|0.0|0.0|1.0|0.0|Jim Cramer: Boeing tweet confirms trump as negotiator-in - USA TODAY https://t.co/gnyTLFSkHH
testrssnews|bbc|0.0|0.0|1.0|0.0|Trump on Twitter https://t.co/XPBsNQ7pSt
NMatte33|youlivethrice|0.4926|0.0|0.715|0.285|"RT @youlivethrice: We're back, thanks to Trump! #MerryChristmas https://t.co/VltY2nTw7D"
NMatte33|twitter|0.4926|0.0|0.715|0.285|"RT @youlivethrice: We're back, thanks to Trump! #MerryChristmas https://t.co/VltY2nTw7D"
matometrump|trump|0.0|0.0|1.0|0.0|   https://t.co/zouJ8fejYz
PedroCo16889625|kurteichenwald|0.5574|0.0|0.847|0.153|"RT @kurteichenwald: If Trump started getting praise 4  appointments from ISIS, do you think Fox News would start running stories about how"
mharvey816|SeanMcElwee|0.6249|0.0|0.796|0.204|"RT @SeanMcElwee: Trump gave cabinet positions to 6 major donors, which is unprecedented. Great reporting from @mateagold. https://t.co/2w4v"
mharvey816|t|0.6249|0.0|0.796|0.204|"RT @SeanMcElwee: Trump gave cabinet positions to 6 major donors, which is unprecedented. Great reporting from @mateagold. https://t.co/2w4v"
jennifer4nm|kurteichenwald|0.7089|0.0|0.772|0.228|"RT @kurteichenwald: Trump says: So smart doesnt need daily intel briefings, knows more about ISIS than military, knows tax code better than"
cynthia_gail|Suthen_boy|-0.5106|0.155|0.845|0.0|"RT @Suthen_boy: Trump bashes CIA, dismisses Russian hacking report https://t.co/YQCXz2jSA3 He knows what corrupt liar O is pulling #tcot #p"
cynthia_gail|usatoday|-0.5106|0.155|0.845|0.0|"RT @Suthen_boy: Trump bashes CIA, dismisses Russian hacking report https://t.co/YQCXz2jSA3 He knows what corrupt liar O is pulling #tcot #p"
mrmarkplum|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
TheRick35|bfraser747|0.7003|0.0|0.726|0.274|"RT @bfraser747: ""To say that the Russians would like 2 have Trump? Look, the Russians have been playing this administration like a fiddle"""
trump_woman|eggvatar|0.0|0.0|1.0|0.0|@eggvatar John Bolton is NOT in show biz so here's his Bio for your edification. Bolton is SOS Candidate for Trump. https://t.co/NZcdkkGq01
trump_woman|twitter|0.0|0.0|1.0|0.0|@eggvatar John Bolton is NOT in show biz so here's his Bio for your edification. Bolton is SOS Candidate for Trump. https://t.co/NZcdkkGq01
laurenm|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
thePoWer_RangeR|NBCNews|0.7579|0.0|0.698|0.302|"RT @NBCNews: CIA concludes Russia mounted covert operation to help Trump win, congressional official says https://t.co/hHlhMGJgwL https://t"
thePoWer_RangeR|nbcnews|0.7579|0.0|0.698|0.302|"RT @NBCNews: CIA concludes Russia mounted covert operation to help Trump win, congressional official says https://t.co/hHlhMGJgwL https://t"
LisaToddSutton|dwaynecobb|0.7096|0.0|0.781|0.219|RT @dwaynecobb: ....    So Russia gives election to Trump &amp; Russia gets Tillerson at State and Flynn as National Security Adviser as a bonus
JHSaunders|funder|0.0|0.0|1.0|0.0|RT @funder: Breaking:Trump started doing business in Taiwan in 2008 #TrumpLeaks#FridayFeeling #msnbc #cnn @JoyAnnReid @maddow @Lawrence @c
NateInPhilly|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
eNewsPR_DK|b|0.0|0.0|1.0|0.0|Donald Trump varsler opgr med USA's et-Kina-politik https://t.co/rYLsgKYXyA #nyheder #News
Isabel__Jones|RealRussBaker|0.4576|0.0|0.875|0.125|"RT @RealRussBaker: When even CIA and NSA think Trump and his Strangeloves are wacko, you know things are gonna get more interesting"
Web20watch|politico|0.0|0.0|1.0|0.0|Trump blasts NBC on Twitter - Politico https://t.co/yjrZ8ygjie
chuckbrixey|realDonaldTrump|-0.9349|0.461|0.475|0.064|@realDonaldTrump @NBCNightlyNews @CNN shut the fuck up Trump you piece of shit it sucks when they print the truth huh you lying bastard
thegranolamom|MMFlint|-0.4767|0.256|0.744|0.0|@MMFlint youtube riddled with fake comments on trump videos https://t.co/mXOPLfJCmb
thegranolamom|youtube|-0.4767|0.256|0.744|0.0|@MMFlint youtube riddled with fake comments on trump videos https://t.co/mXOPLfJCmb
ramsay_scott|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: Media: ""Trump's racist""""Trump's fascist""""Trump's sexist""""Trump's hitler""""Trump's a clown""""Trump's not serious"""""
TurnTNBlue|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: Trump: 'Nobody really knows' if #ClimateChange is real. Um... Apart from every scientist who works on the subject?! Idi
LKuehn4|kurteichenwald|0.126|0.146|0.687|0.167|"RT @kurteichenwald: Putin staff consultant re: Trump choices: ""This is a fantastic team!""Remember when Romney said Russia biggest threat?"
pisannd5|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: When Obama used Dijon mustard, Fox attackd him 4 not using yellow mustrd (true) Yet they shrug when Trump says doesnt n"
pulpmarkets|bloomberg|-0.34|0.156|0.844|0.0|markets: RT business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/nKcrVkG16N https://t.co/97oXvEhFa9
Dewblue1|TheDonaldNews|0.128|0.111|0.754|0.136|RT @TheDonaldNews: FBI Investigation Refutes CIA=&gt; Theres No Evidence Russia Tried to Help Trump https://t.co/lUPBb1wd0y #FoxNews #Tucker
Dewblue1|thegatewaypundit|0.128|0.111|0.754|0.136|RT @TheDonaldNews: FBI Investigation Refutes CIA=&gt; Theres No Evidence Russia Tried to Help Trump https://t.co/lUPBb1wd0y #FoxNews #Tucker
Adriene26|AriMelber|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
Adriene26|t|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
ibleedandstuff|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
RWNemanich|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
SkyLaser3|abctweet100|-0.7845|0.345|0.655|0.0|RT @abctweet100: Trump's Antagonistic Rhetoric Towards China is Dangerous-His Lack of Diplomacy Shows Inexperience &amp; Stupidity #News  https
plowman_robert|CarlBullock16|-0.5574|0.194|0.806|0.0|RT @CarlBullock16: Trump-Themed Star Wars Posters Featuring MILO Spotted Around Rogue One Premiere Area https://t.co/B34ZMfBMLX https://t
plowman_robert|breitbart|-0.5574|0.194|0.806|0.0|RT @CarlBullock16: Trump-Themed Star Wars Posters Featuring MILO Spotted Around Rogue One Premiere Area https://t.co/B34ZMfBMLX https://t
Synergism3|JuddLegum|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
Synergism3|t|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
thisischrisb|voxdotcom|-0.3252|0.163|0.837|0.0|Donald Trump is running the least popular transition in decades https://t.co/PQcc5AoQjL via @voxdotcom
thisischrisb|vox|-0.3252|0.163|0.837|0.0|Donald Trump is running the least popular transition in decades https://t.co/PQcc5AoQjL via @voxdotcom
LibbySwenson|swin24|-0.0572|0.055|0.945|0.0|"RT @swin24: Today, Trump says he doesnt want anyone hacking the U.S.In July, he called on Russia to hack the U.S. govt.https://t.co/"
EricBryan7|YouTube|0.3182|0.0|0.859|0.141|The Real Truth Behind The CIA Report Of Russian Hacking Electing Trump https://t.co/9BQBMwGGmP via @YouTube
EricBryan7|youtube|0.3182|0.0|0.859|0.141|The Real Truth Behind The CIA Report Of Russian Hacking Electing Trump https://t.co/9BQBMwGGmP via @YouTube
bbdevices|tribelaw|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
bbdevices|twitter|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
inklake|EricBoehlert|0.0|0.0|1.0|0.0|RT @EricBoehlert: Trump can't find a single senior intel official to step forward and say Russia absolutely not involved in election?
INSOMNIAK_DJ|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
NetaniaLim|davidfolkenflik|0.0|0.0|1.0|0.0|RT @davidfolkenflik: Did not expect this exegesis of gaslighting and its relationship to current day politics from Teen Vogue https://t.co/
NetaniaLim|t|0.0|0.0|1.0|0.0|RT @davidfolkenflik: Did not expect this exegesis of gaslighting and its relationship to current day politics from Teen Vogue https://t.co/
llostgirl|ghefrentte|0.0|0.0|1.0|0.0|RT @ghefrentte: Quando tem brasileiro apoiando o Trump na timeline https://t.co/PzmbxQaAhb
llostgirl|twitter|0.0|0.0|1.0|0.0|RT @ghefrentte: Quando tem brasileiro apoiando o Trump na timeline https://t.co/PzmbxQaAhb
ArmstrongLance3|elijahdaniel|0.7579|0.0|0.683|0.317|RT @elijahdaniel: that time I became a best selling author because I wrote a 20 page trump erotic novel https://t.co/DSq421WtkJ
ArmstrongLance3|twitter|0.7579|0.0|0.683|0.317|RT @elijahdaniel: that time I became a best selling author because I wrote a 20 page trump erotic novel https://t.co/DSq421WtkJ
rolmarjr|mobile|0.4767|0.0|0.846|0.154|The Washington Post and The New York Times reported on Friday that American intelligence agencies had concluded... https://t.co/T1VSGIBRjQ
innaroz|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
gooberspa|Nate_Cohn|0.1531|0.121|0.738|0.141|RT @Nate_Cohn: I guess the Trump-Bolton case is that there were 2m illegal votes and a CIA false flag op in one of the greatest victories i
themayorofoc|V_of_Europe|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
themayorofoc|thegatewaypundit|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
agscribbler|TheRickWilson|0.0|0.0|1.0|0.0|"RT @TheRickWilson: The word ""intelligence"" doesn't mean what Donald Trump thinks it means in this case https://t.co/Nxsmr3770D"
agscribbler|time|0.0|0.0|1.0|0.0|"RT @TheRickWilson: The word ""intelligence"" doesn't mean what Donald Trump thinks it means in this case https://t.co/Nxsmr3770D"
ScienceWorld9|itechpost|0.0772|0.0|0.894|0.106|What Future Awaits The Science Department Under Trump Administration? - iTech Post https://t.co/n7AuypEgSY
DiMill46|paulkrugman|0.7269|0.0|0.757|0.243|"RT @paulkrugman: Between Comey and the popular vote, you can make a strong case that Trump victory was fundamentally illegitimate. But wher"
lobster_dog|thesilentshore|0.0|0.0|1.0|0.0|@thesilentshore someone from Trump's campaign has it
TaiwanNewsshow|nytimes|0.0|0.0|1.0|0.0|Trump Suggests Using Bedrock China Policy as Bargaining Chip - New York Times https://t.co/xXMYtBPAjI
worldnews134|bbc|0.0|0.0|1.0|0.0|Trump on Twitter https://t.co/tDs5YV8EXt
DessyFenix|ericgarland|0.6059|0.075|0.746|0.179|"RT @ericgarland: Trump - a moron - is probably unlikely to take the whole enchilada, but that's perfect. If he gets close enough, he can cr"
DespinaKaddouri|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
GlennLittle5|dmartosko|0.0|0.0|1.0|0.0|RT @dmartosko: DOCUMENTS: Trump was RIGHT about $4+ billion cost for new Air Force One planes https://t.co/TaHdJGufsN via @MailOnline
GlennLittle5|dailymail|0.0|0.0|1.0|0.0|RT @dmartosko: DOCUMENTS: Trump was RIGHT about $4+ billion cost for new Air Force One planes https://t.co/TaHdJGufsN via @MailOnline
respectinc|jayrosen_nyu|-0.3182|0.121|0.879|0.0|RT @jayrosen_nyu: 5/ From Trump a steady flow of easy-to-check lies as both a show of power and to cast the press in the role of petty but
NicoleCynLane|ananavarro|-0.1027|0.136|0.746|0.118|"RT @ananavarro: Been off-line for hours vicariously suffering @MiamiDolphins' game...tell me, has Trump named Putin ""Special Advisor to the"
cbrownx|mikandynothem|0.3802|0.088|0.767|0.146|RT @mikandynothem: Ruth Bader Ginsburg said she would resign if Trump won. Hit the road lady! That will give Trump even more Conservatives
ckensingtn|AriFleischer|-0.7351|0.212|0.788|0.0|"RT @AriFleischer: If it's wrong for Trump 2receive royalties as EP of his TV show, was it wrong for Obama and Hillary 2receive royalties fo"
yytirado|Reuters|0.0|0.0|1.0|0.0|RT @Reuters: McCain to Trump on Russian hacking: 'The facts are there' - CBS https://t.co/QoesspVeoq https://t.co/pP6xj54U5Q
yytirado|reuters|0.0|0.0|1.0|0.0|RT @Reuters: McCain to Trump on Russian hacking: 'The facts are there' - CBS https://t.co/QoesspVeoq https://t.co/pP6xj54U5Q
knew777771|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
knew777771|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
Hehe24Small|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
walkileaks|newsyarn|0.0|0.0|1.0|0.0|"Despite scientific consensus, Trump says nobody knows if climate change isreal https://t.co/JmMs384wfv"
Dina_Tan73|FieldDiamond|0.3612|0.0|0.865|0.135|@FieldDiamond @TheBudgetGuy @RuthMarcus we'll never know with a malignant narcissist and a sociopath like Trump ppl are disposable 4 him
alfredenmn|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
FaithFlaherty3|jmaboshie|0.8573|0.165|0.482|0.354|"RT @jmaboshie: Im Vladimir, i stole the election for #Trump but I let Hillary win the popular vote. I forgot to rig that part. My bad. Won'"
Anj_T|liamstack|0.0772|0.105|0.739|0.156|RT @liamstack: Now that Twitter has cracked down on the pro-Trump bots the top replies to @realDonaldTrump are mostly comedians mocking him
laurine3215|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
tammy_wesa|DavidCornDC|0.0|0.0|1.0|0.0|RT @DavidCornDC: Why Donald Trump appointing John Bolton to any post is crazy...even for Trump: https://t.co/KjbZP4B4Z3
tammy_wesa|m|0.0|0.0|1.0|0.0|RT @DavidCornDC: Why Donald Trump appointing John Bolton to any post is crazy...even for Trump: https://t.co/KjbZP4B4Z3
rachmanworks|CNBC|0.0|0.0|1.0|0.0|RT @CNBC: BREAKING: Trump picks Exxon Mobil CEO Tillerson to be his Secretary of State - @NBCNews
OnlineMarketmix|politico|0.0|0.0|1.0|0.0|Trump blasts NBC on Twitter - Politico https://t.co/QT0I53g8RT
HelenEckard|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
mindburnr|AdamVanBavel|0.169|0.115|0.733|0.152|"RT @AdamVanBavel: Trump doesn't need security briefings because he's 'like, a smart person'  #DumpTrump #YoureFired https://t.co/NkuAO9xfI"
mindburnr|t|0.169|0.115|0.733|0.152|"RT @AdamVanBavel: Trump doesn't need security briefings because he's 'like, a smart person'  #DumpTrump #YoureFired https://t.co/NkuAO9xfI"
mzbitca|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
mzbitca|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
Habanera119|Bipartisan|-0.2808|0.18|0.695|0.124|"BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/XfHyZsE7bf via @Bipartisan Report"
Habanera119|bipartisanreport|-0.2808|0.18|0.695|0.124|"BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/XfHyZsE7bf via @Bipartisan Report"
cookiebucky1|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
cookiebucky1||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
Zwelkiss|helenmaryme|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
Zwelkiss|twitter|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
MaelinnHughes|tomtomorrow|-0.7841|0.247|0.703|0.05|RT @tomtomorrow: Thought of what Trump's election means for this country has left me feeling the sort of grief I have felt after death of s
asbinvancity|PattyParsonsPat|0.0|0.0|1.0|0.0|RT @PattyParsonsPat: Lmbo my tweet seen by more people than Donald trump got votes https://t.co/gChAKEjEKh
asbinvancity|twitter|0.0|0.0|1.0|0.0|RT @PattyParsonsPat: Lmbo my tweet seen by more people than Donald trump got votes https://t.co/gChAKEjEKh
HURRICANEPAUL|stranahan|0.7506|0.0|0.701|0.299|".@stranahan These ""rebels"" are going to wish Hillary won after President Trump is finished with them.#WalkingDead @YouTube"
EnvironmenLaw|politico|0.0|0.0|1.0|0.0|"'I'm very open-minded on environment,' Trump says - Politico https://t.co/oRBSjNto0W"
FactsVsOpinion|ginammack|0.0|0.0|1.0|0.0|RT @ginammack: @Bencjacobs And it's just coincidence that the Trump cabinet is pro-Russia?
SOS_1313|mitchellvii|0.7914|0.108|0.56|0.332|"RT @mitchellvii: I would not be surprised if Russia favored Trump winning.  After 8 years, they didn't want another idiot running America."
trumpsquatch|trumpsquatch|0.0|0.0|1.0|0.0|RT @trumpsquatch: Boomsticks for trump #MAGA #2A @girlswithguns_ @HotGirlsAndGuns #guns #bikini https://t.co/TS1rPWCbEu
trumpsquatch|twitter|0.0|0.0|1.0|0.0|RT @trumpsquatch: Boomsticks for trump #MAGA #2A @girlswithguns_ @HotGirlsAndGuns #guns #bikini https://t.co/TS1rPWCbEu
zweckfam|LOLGOP|-0.6917|0.248|0.67|0.082|RT @LOLGOP: Trump doesn't like to be known as the biggest popular vote loser to be elected in modern history. It would be rude to point tha
RebelHeartWorld|StopTrump2020|0.0|0.0|1.0|0.0|"RT @StopTrump2020: #Trump filling his cabinet with #FriendsOfPutin, UNQUALIFIED swamp creatures, Billionaires and big donors.  #NotMyPresid"
PTsully55|cutasterfee|0.0|0.0|1.0|0.0|@cutasterfee for mother Russia.. your a trump agent
GarronRobert|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
GarronRobert|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
DhitaPuss|punyakitasemuanih|0.0|0.0|1.0|0.0|" https://t.co/jowkYMygu3  #bokep #bispak Baru  Info Baca Melania Trump Blak-blakan Soal Ranjang, Ternyata Begini Donald Trump di Atas "
snarkysyntax|meganamram|0.0|0.0|1.0|0.0|RT @meganamram: Real question: does Trump believe in object permanence
Nuwanda9|KeepAmerGr8|-0.4939|0.167|0.833|0.0|RT @KeepAmerGr8: Trump Thinks Daily Briefings Are For Losersand Other Scary Revelations About His Management Philosophy https://t.co/hlj9H
Nuwanda9|t|-0.4939|0.167|0.833|0.0|RT @KeepAmerGr8: Trump Thinks Daily Briefings Are For Losersand Other Scary Revelations About His Management Philosophy https://t.co/hlj9H
Bayathread|msfoundation|0.5859|0.0|0.703|0.297|@msfoundation follow @RachelleHodgs for brilliant graphing of Trump word salads.
NikkiNiceOKC|AP|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
NikkiNiceOKC|t|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
debesponomi|HamiltonElector|-0.4401|0.115|0.843|0.042|RT @HamiltonElector: RT The only thing that matters now is educating EVERYONE that Donald Trump is not President yet. He has not won. #Dec1
AZULCAMPEON10|politicomx|0.0|0.0|1.0|0.0|"RT @politicomx: #Trump se declar ""gran creyente"" del libre comercio. Por lo mismo, gravar a las empresas que salgan de #EUA: https://t.c"
AZULCAMPEON10||0.0|0.0|1.0|0.0|"RT @politicomx: #Trump se declar ""gran creyente"" del libre comercio. Por lo mismo, gravar a las empresas que salgan de #EUA: https://t.c"
DeDimacrow|politico|0.5893|0.0|0.797|0.203|"This is the Soft ball BS LOL Not news from Fox,the BS Not new network! https://t.co/9TH8qDW0lT"
downtown7thave|Toure|0.6647|0.113|0.532|0.355|RT @Toure: Trump says he doesnt need intelligence briefings because Im a smart person. God save us.
ceili_woman|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
mtighe15|USARedOrchestra|-0.836|0.294|0.706|0.0|"RT @USARedOrchestra: When u equate emails w/ racism, misogyny, sexual assault &amp; 10x more coverage than any single trump story, then check s"
notjustwarri|twitter|-0.2732|0.139|0.861|0.0|"#notjustwarriPolitics|Trump's Expected Labor Pick, Andrew Puzder, Is Minimum Wage Critic - New York Times https://t.co/9ulaBeQOec"
JoeFeagin|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
JoeFeagin|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
Rene_Berto|amazon|0.0|0.0|1.0|0.0|Trump aegri somnia beati possidentes #linenews #holidayswithheart https://t.co/DG7SwspZTX https://t.co/5EyCSScuSN
jayawells|calatayud7|0.0|0.0|1.0|0.0|RT @calatayud7: We cannot let this go.  The future of America is at stake.  Trump cannot take office. https://t.co/L9ySOQNc8O
jayawells|twitter|0.0|0.0|1.0|0.0|RT @calatayud7: We cannot let this go.  The future of America is at stake.  Trump cannot take office. https://t.co/L9ySOQNc8O
Melanymlove|nytimes|-0.296|0.285|0.57|0.146|"Abortion Foes, Emboldened by Trump, Promise Onslaught of Tough Restrictions https://t.co/GZ9XuRNT87 https://t.co/5gOm2ykgDr"
retrotimewarp|SamGrittner|0.0|0.0|1.0|0.0|@SamGrittner Yet another potential  whack job choice for the Trump cabal.
Egy_U|nytimes|0.0|0.0|1.0|0.0|"Boeing Seeks to Sell Planes to Iran, and the Deal to Trump https://t.co/v6blCUDDlc"
SeriesaddictIra|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Bitch_Wear|Ali_Tmak_Store.https//t.co/qLTFpnmhtt|0.0|0.0|1.0|0.0|............ President Trump tShirts...................... by Ali Tmak------------&gt; @Ali_Tmak_Store.https://t.co/qLTFpnmhtt
seanskiwords|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
TechNewsDB|technewsdb|0.0|0.0|1.0|0.0|"Larry Page, Tim Cook said to attend Donald Trump's tech summit     - CNET - https://t.co/DtABAjRNS0 https://t.co/MaoLhXLySG"
PatPatojson|Corporatocrazy|-0.765|0.32|0.68|0.0|RT @Corporatocrazy: Lunatic Loser Liberals trying to stage a coup by using Russia conspiracy#Trump #CIA #FBI https://t.co/WEcIzKtb8X
PatPatojson|naturalnews|-0.765|0.32|0.68|0.0|RT @Corporatocrazy: Lunatic Loser Liberals trying to stage a coup by using Russia conspiracy#Trump #CIA #FBI https://t.co/WEcIzKtb8X
lynndals|CaptainsLog2016|-0.5423|0.276|0.623|0.101|"RT @CaptainsLog2016: Dear @CanadaCan I book a 4 year stay in your country?I have no felonies, I pay taxes, and I didn't vote for Trump"
JoeRash3|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
JoeRash3|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
danaarsenault|twitter|0.0|0.0|1.0|0.0|RIP Patriotic Pepe. AKA the Russian bot who commented first under every Trump tweet for over a year. https://t.co/FgJDUshtGj
USSenateview|thehill|-0.3875|0.193|0.807|0.0|Dem senator to Trump: Russia is not our friend - The Hill https://t.co/svNantc7zK
Floridaartist1|SandraTXAS|0.8126|0.0|0.549|0.451|RT @SandraTXAS: Trump loves AmericaObama loves communism and dictators #MAGA#AmericaFirst#WeekendUpdate https://t.co/nt6SBJL9Bf
Floridaartist1|twitter|0.8126|0.0|0.549|0.451|RT @SandraTXAS: Trump loves AmericaObama loves communism and dictators #MAGA#AmericaFirst#WeekendUpdate https://t.co/nt6SBJL9Bf
madelineloveg|nytimes|-0.296|0.285|0.57|0.146|"Abortion Foes, Emboldened by Trump, Promise Onslaught of Tough Restrictions https://t.co/g3D2u7m56j https://t.co/QUUCzd4WyS"
iPhonefanclubs|appleinsider|0.0|0.0|1.0|0.0|Apple's Tim Cook among tech executives meeting with Donald Trump on Wednesday - report - AppleInsider (press https://t.co/SaPPITR4Hh
mcmisher|GeorgeTakei|-0.1779|0.182|0.694|0.123|"RT @GeorgeTakei: The Russians hacked the RNC but didn't release those emails. They wanted to help Trump get elected, but could threaten him"
LibraQueenLibby|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
LibraQueenLibby|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
DebbiebB15|VampKiraLynn|-0.4215|0.144|0.778|0.078|RT @VampKiraLynn: @funder @kellyannepolls America as we know it will die the day trump takes the office. This will NOT end well. #Resist
ramaiamar|yahoo|-0.0772|0.098|0.902|0.0|Three Decades Of Trump's Russian Ties Exposed In One Democratic Coalition Report https://t.co/B0ciyj1sKl
padilloh|ebromleymdphd|0.4389|0.0|0.804|0.196|"RT @ebromleymdphd: @jayrosen_nyu yes, I agree! at first, I didn't quite get it but I keep returning to it. from: https://t.co/jplWaAccJ7"
padilloh|qz|0.4389|0.0|0.804|0.196|"RT @ebromleymdphd: @jayrosen_nyu yes, I agree! at first, I didn't quite get it but I keep returning to it. from: https://t.co/jplWaAccJ7"
PeterTownsend7|ptbooks|0.5106|0.0|0.752|0.248|The 'Prophet' and Free Speech  #trump #maga #isis #pjnet https://t.co/zAhdl485xH https://t.co/yenXR9Duus
corytheswirler|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
SmarterThanAl1|smarterthanalbert|0.4515|0.0|0.815|0.185|What are your thoughts on elected President #Trump? Will he keep his promises? https://t.co/GgkZgFzgNq
GuruMarketeer|smarterthanalbert|0.4515|0.0|0.815|0.185|What are your thoughts on elected President #Trump? Will he keep his promises? https://t.co/fZdbDFUe1N
RNRoxx|HamiltonElector|0.2298|0.123|0.757|0.12|"RT @HamiltonElector: Mr. Trump you are hardly a genius, no matter what Comrade Putin says.  We are smarter than you. We are #hamiltonelecto"
Pixelfish|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
thebitterfig|JoyAnnReid|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
thebitterfig|twitter|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
TrumpNation10|Sammie_Snickers|-0.296|0.167|0.833|0.0|RT @Sammie_Snickers: Trump's Pennsylvania Electors Showing No Signs Of Flipping https://t.co/YVU403TFe0@mitchellvii @gatewaypundit
TrumpNation10|philadelphia|-0.296|0.167|0.833|0.0|RT @Sammie_Snickers: Trump's Pennsylvania Electors Showing No Signs Of Flipping https://t.co/YVU403TFe0@mitchellvii @gatewaypundit
captainolya|janiobi|-0.6428|0.2|0.8|0.0|"RT @janiobi: Oh man this shit about Casey Affleck. I mean, Nate Parker. I mean, President Elect Donald Trump. I mean..."
jane_spillane|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
cvasilevski|Evan_McMullin|0.0119|0.094|0.81|0.096|RT @Evan_McMullin: It must be clear that Donald Trump is not a loyal American and we should prepare for the next four years accordingly. @r
Scrutinator|andres20ad|-0.296|0.104|0.896|0.0|"@andres20ad @OdetteEngel Ms tolerancia, amigo. Si Trump gan en democracia, donde gana la mayora y no las minoras, TODO es posible."
OKCliberal|nbcnews|0.7579|0.0|0.606|0.394|"Russia mounted a covert operation to help Trump win, source tells NBC https://t.co/3XFwvO4RL4"
grannyso|melreynoldsU|-0.5927|0.129|0.871|0.0|RT @melreynoldsU: Your ego won't let you Trump but pull this Exxon guy. It will be your first major embarrassment if you put him up for Sec
ballerinaX|leahmcelrath|0.0|0.0|1.0|0.0|"RT @leahmcelrath: This is a thorough compilation on @dailykos of resources regarding Putin, Dugin, Spencer, Bannon, and Trump:https://t.c"
ballerinaX||0.0|0.0|1.0|0.0|"RT @leahmcelrath: This is a thorough compilation on @dailykos of resources regarding Putin, Dugin, Spencer, Bannon, and Trump:https://t.c"
yoenterado|youtube|0.0|0.0|1.0|0.0|Los mejores memes del debate Clinton vs Trump https://t.co/O7sioTluO4  #FelizDomingo
scott_boore|twitter|-0.2411|0.164|0.836|0.0|Trump wouldn't know truth if it hit in the face. https://t.co/TBhKmNjMuL
donkrusty|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
nancy73gg|amrightnow|0.0|0.0|1.0|0.0|"RT @amrightnow: Big big wall"" Make Video #1 (Trump About You) https://t.co/j58e8aacrE #WisconsinPrimary #Wisconsin #Wisconsinpoll https://t"
nancy73gg|youtube|0.0|0.0|1.0|0.0|"RT @amrightnow: Big big wall"" Make Video #1 (Trump About You) https://t.co/j58e8aacrE #WisconsinPrimary #Wisconsin #Wisconsinpoll https://t"
lisatalley045|asamjulian|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
lisatalley045|twitter|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
DermArch|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
DermArch||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
AngelicPrado|LightsOut2017|-0.2732|0.129|0.796|0.075|"RT @LightsOut2017: Exclusive: Billionaire green activist Steyer vows to battle Trump, says money not an issue https://t.co/EncAeeZuUw via @"
AngelicPrado|reuters|-0.2732|0.129|0.796|0.075|"RT @LightsOut2017: Exclusive: Billionaire green activist Steyer vows to battle Trump, says money not an issue https://t.co/EncAeeZuUw via @"
MLBDenver|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
MLBDenver||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
gkilday|ABFalecbaldwin|0.886|0.059|0.472|0.469|Uh-0h. @ABFalecbaldwin just won a CritcsChoice Award for playing Trump. Hope @realDonaldTrump isn't watching or he'll demand a recount
erinhale|dpa_intl|0.0|0.0|1.0|0.0|RT @dpa_intl: US president-elect Donald Trump in an interview with Fox News defends his decision to select several retired generals for his
yuweile|wikileaks|-0.296|0.091|0.909|0.0|RT @wikileaks: No link between Trump &amp; RussiaNo link between Assange &amp; RussiaBut Podesta &amp; Clinton involved in selling 20% of US uranium
miscelaineee|KeithOlbermann|0.0|0.0|1.0|0.0|RT @KeithOlbermann: CIA revealed Russia HAD tampered for Trump. From 10/14: when Trump revealed he knew HOW they were doing it for him http
yardsailor43|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
Lisa_Iannucci|JohnFPfaff|-0.0516|0.095|0.905|0.0|"RT @JohnFPfaff: So if each daily briefing says ""Russians are ten miles closer to Warsaw than yesterday,"" how long after Warsaw falls will T"
vdutat|HamiltonElector|-0.4401|0.115|0.843|0.042|RT @HamiltonElector: RT The only thing that matters now is educating EVERYONE that Donald Trump is not President yet. He has not won. #Dec1
DessyFenix|ericgarland|-0.529|0.189|0.811|0.0|RT @ericgarland: The Russians didn't create Trump - only New York City and American gullibility could have done that.But they've got a SW
robertmeyer9|socialmaze|-0.5994|0.245|0.755|0.0|Cultural War and the Election of Donald Trump  https://t.co/upeJYLKbhQ  #conservatives #liberals #progressives https://t.co/3MRkf9gCru
Reforma|reforma|-0.34|0.13|0.87|0.0|La comunidad de inteligencia de EU se alarm ante los comentarios y el rechazo de Donald Trump https://t.co/KkzGp0BLjt
caroljdavy|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
kayewhitehead|kayewisewhitehead|-0.1027|0.167|0.833|0.0|"Trump and Gender Bias, By theNumbers https://t.co/zaTRbRVvuK https://t.co/yxXVrUMiqq"
furngals2|DailyCaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
furngals2|dailycaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
gaga20219gs|amjoyshow|0.0|0.0|1.0|0.0|RT @amjoyshow: Scott Dworkin (@FUNDER) joins on #TrumpLeaks &amp; #DworkinReport that consolidates all Donald Trump's Russian ties over many ye
BenReclused|StoneColdTruth|0.4404|0.099|0.673|0.229|"RT @StoneColdTruth: https://t.co/mnsZmkBMN9Corprations around the country claim there is no local talent, that they NEED H1-B. Pray tell,"
BenReclused|t|0.4404|0.099|0.673|0.229|"RT @StoneColdTruth: https://t.co/mnsZmkBMN9Corprations around the country claim there is no local talent, that they NEED H1-B. Pray tell,"
angulosiete|angulo7|0.0|0.0|1.0|0.0|#Economa #Canaive abrir oficina en #EU pese a poltica antimigratoria de #Trump | ngulo 7 https://t.co/tgmastUnh9
THE_DAILY_BLEAT|DailyCaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
THE_DAILY_BLEAT|dailycaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
mdjtraveler|KellyannePolls|0.6808|0.0|0.763|0.237|@KellyannePolls @AmerPride777 Lil' Marco &amp; stooges better get in line or face the Trump wrath. Trump's voters support Trump @realDonaldTrump
rockshout|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
catoletters|veteranstoday|-0.5719|0.316|0.684|0.0|2015 McCain's Treasonous Can of Worms via https://t.co/uSxnxp7IRH:  https://t.co/0hrGMk1kqQ
lehudgins|MattOrtega|0.0|0.0|1.0|0.0|Corrupt AF: 12 hours since the latest report of corruption by Donald Trump. https://t.co/XFeTmsISeF via @MattOrtega
lehudgins|corrupt|0.0|0.0|1.0|0.0|Corrupt AF: 12 hours since the latest report of corruption by Donald Trump. https://t.co/XFeTmsISeF via @MattOrtega
RevPastorJack|ijr|0.0|0.0|1.0|0.0|Time to overhaul the CIA and other government offices. https://t.co/zOX6kaNljq
ConservativLuke|unsavoryagents|0.0|0.0|1.0|0.0|RT @unsavoryagents: PREPARE FOR THE LEFT TO TAKE A COLLECTIVE SHIT!!!https://t.co/WuQaHWBhsq
ConservativLuke|nbcnews|0.0|0.0|1.0|0.0|RT @unsavoryagents: PREPARE FOR THE LEFT TO TAKE A COLLECTIVE SHIT!!!https://t.co/WuQaHWBhsq
holtmapa|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
holtmapa||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
openomroep|nbcnews|-0.4939|0.325|0.515|0.16|#news Intelligence Agencies Distressed by Trump's Rejection of Findings on Russia - NBCNews https://t.co/vRmEF45Tvz
MickBlair54|breitbart|-0.34|0.156|0.844|0.0|Gavin Newsom: Trump's Election a 'Leap Backward' for States with Stringent Gun Control - Breitbart https://t.co/6oYoQISc9n
amcnair00|nbcnews|0.0|0.0|1.0|0.0|https://t.co/Kb8ExVre86
blueinthesouth|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
Phil_Laird1|VoteHillary2016|0.0|0.0|1.0|0.0|"RT @VoteHillary2016: Trump's Secretary of State pick, @Exxon's @rex_tillerson, toasting Putin &amp; associates after signing lucrative deal. ht"
addykateglen|ReaganBattalion|-0.5719|0.281|0.719|0.0|"RT @ReaganBattalion: .@oreillyfactor accused @GeorgeWill in ""undermining conservatism"" for opposing Trump. @JudgeJeanine: Opposing Trump"
lonegamer78|benschwartzy|-0.5177|0.218|0.66|0.122|"RT @benschwartzy: It only took one FBI agent to ruin Nixon (Felt) and one to ruin Hillary (Comey). So, I'm very happy to see Trump making a"
sasachio72|tackettdc|0.296|0.0|0.896|0.104|"RT @tackettdc: ""Russia, they said, had intervened with the primary aim of helping make Donald J. Trump president"" @markmazzettinyt  https:/"
sasachio72||0.296|0.0|0.896|0.104|"RT @tackettdc: ""Russia, they said, had intervened with the primary aim of helping make Donald J. Trump president"" @markmazzettinyt  https:/"
burghline|burghline|0.4215|0.0|0.823|0.177|Netanyahu says he hopes to work with Trump to undo Iran deal https://t.co/NJm6rlA9J6 https://t.co/esvxaDXvwL
anobscureartist|TheEconomist|0.34|0.119|0.693|0.188|"RT @TheEconomist: Republicans are denying that Russias authoritarian, anti-American government wanted Mr Trump to win https://t.co/WGgzEMk"
anobscureartist|t|0.34|0.119|0.693|0.188|"RT @TheEconomist: Republicans are denying that Russias authoritarian, anti-American government wanted Mr Trump to win https://t.co/WGgzEMk"
IntrovertRN1975|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
IntrovertRN1975|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
Deplorablefrog1|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
ZeliaLH|BV|-0.1926|0.118|0.8|0.082|"#Chinese investors aren't flustered by #Trumpophobia; esp., when they are the biggest holders of #US debt https://t.co/HqiApX6TII via @BV"
ZeliaLH|linkis|-0.1926|0.118|0.8|0.082|"#Chinese investors aren't flustered by #Trumpophobia; esp., when they are the biggest holders of #US debt https://t.co/HqiApX6TII via @BV"
crownlifelive|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
GREEN_THE_WORLD|m|0.0|0.0|1.0|0.0|Trump confirme son scepticisme concernant le changement climatique - 7sur7 https://t.co/ii30EcP2Ml
lollytw|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
lollytw|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
imagin8ion|behindyourback|0.5423|0.088|0.696|0.216|"RT @behindyourback: Look, Trump's just too busy to bother with intelligence briefings on the fundamental safety of our country and its citi"
Quietness_Trust|MrJonCryer|-0.4019|0.114|0.886|0.0|"RT @MrJonCryer: And for those Trump Voters who thought there was something nefarious about Hillary's emails, why are you ignoring all this?"
vincicat|tomphillipsin|-0.7783|0.264|0.736|0.0|"RT @tomphillipsin: Beijing life, late 2016: wake up, inhale smog, think, 'What the hell did Donald Trump say while I was sleeping?'"
Shanny_resqchi|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
PatriotJane2|davidfrum|-0.4019|0.186|0.722|0.093|"@davidfrum Once the Trump admin is in place, they can put political pressure on the special prosecution to make the facts go their way."
emptypockets57|ThePatriot143|0.4466|0.0|0.836|0.164|RT @ThePatriot143: Traitors John McCain and Lindsey Graham JOIN DEMOCRATS to DELEGITIMIZE President-Elect Trump  TruthFeed https://t.co/ne
emptypockets57|t|0.4466|0.0|0.836|0.164|RT @ThePatriot143: Traitors John McCain and Lindsey Graham JOIN DEMOCRATS to DELEGITIMIZE President-Elect Trump  TruthFeed https://t.co/ne
longrunweareall|RadioFreeTom|0.7184|0.0|0.5|0.5|RT @RadioFreeTom: President-elect Trump appreciated your support https://t.co/38ZQbEiaRW
longrunweareall|twitter|0.7184|0.0|0.5|0.5|RT @RadioFreeTom: President-elect Trump appreciated your support https://t.co/38ZQbEiaRW
Damey07|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
melindacasino|mgd4161|-0.0314|0.121|0.765|0.115|RT @mgd4161: @Jamie4Hillary @bluedgal @VABVOX @BernieSanders also played a roll in Trump being elected. I really am not interested n anythi
koalaqueen53|NewYorker|0.0|0.0|1.0|0.0|"RT @NewYorker: If the man who ghostwrote Trump's ""The Art of the Deal"" wrote the book today, he'd call it ""The Sociopath"" https://t.co/tUsH"
koalaqueen53|t|0.0|0.0|1.0|0.0|"RT @NewYorker: If the man who ghostwrote Trump's ""The Art of the Deal"" wrote the book today, he'd call it ""The Sociopath"" https://t.co/tUsH"
CailleachSila|ericgarland|-0.2052|0.114|0.805|0.08|"RT @ericgarland: And now, it's December 11th. Trump says he don't need no stinkin' intel agencies. Russia (BWA HAHAHAHAAAA) blames Ukrain"
Helena83852000|MaxAbrahms|0.0|0.0|1.0|0.0|"RT @MaxAbrahms: Officials familiar with briefings given to Congress say CIA assessment ""wasn't as definitive as has been portrayed."" https:"
NMatte33|SLandinSoCal|-0.7256|0.347|0.481|0.172|"RT @SLandinSoCal: MSNBC caught reporting ""Fake News""! Lying about Trump &amp; Fox. Forced to apologize ON AIR! HaHaHa https://t.co/d6fqf0SkuF"
NMatte33|twitter|-0.7256|0.347|0.481|0.172|"RT @SLandinSoCal: MSNBC caught reporting ""Fake News""! Lying about Trump &amp; Fox. Forced to apologize ON AIR! HaHaHa https://t.co/d6fqf0SkuF"
algegra|huffingtonpost|0.1531|0.16|0.641|0.199|Donald Trump Used To Complain About Obama Not Getting Intelligence Briefings https://t.co/dc2Fteykxg
Maquiavelo61|GobernantesVer|0.0|0.0|1.0|0.0|"Salida de capitales, triunfo de Trump, lento crecimiento y endeudamiento han propiciado vo... https://t.co/MNwFtbFtCp va @GobernantesVer"
Maquiavelo61|gobernantes|0.0|0.0|1.0|0.0|"Salida de capitales, triunfo de Trump, lento crecimiento y endeudamiento han propiciado vo... https://t.co/MNwFtbFtCp va @GobernantesVer"
bbc_fanxyU|nath_celeste|0.0|0.0|1.0|0.0| @nath_celeste  @Nintama_luck  @Prophet_Levi  @mirang_owner @Today_Fortune @Trump_BJ @CSTLT_Fortune
hawaiianlove68|HamiltonElector|0.296|0.083|0.783|0.135|RT @HamiltonElector: Donald Trump trusts InfoWars more than the CIA - let that sink in. He must be stopped #CountryB4Party #CzarNotPOTUS  h
jakerocksalot16|BettyBowers|-0.8309|0.335|0.607|0.057|RT @BettyBowers: TRUMP: Russia hacked DNC. I invite them to hack even more!CIA: Russia hacked even more.TRUMP: The CIA is lying! Russia w
sud_vijay|Redpainter1|0.7703|0.0|0.75|0.25|RT @Redpainter1: Who do you trust: An agency of highly trained intelligence professionals or a man who gets his news from Infowars? https:/
sud_vijay||0.7703|0.0|0.75|0.25|RT @Redpainter1: Who do you trust: An agency of highly trained intelligence professionals or a man who gets his news from Infowars? https:/
stacyllw|twitter|-0.296|0.109|0.891|0.0|"Putin has more knowledge of subversion, espionage, manipulation in his pinky than Trump could ever possess in his e https://t.co/injrSU4A27"
slmbs9|Humans_vs_Trump|-0.2263|0.129|0.783|0.088|"RT @Humans_vs_Trump: Media currently surprised Trump denies Russia hacking.Um, remember when he invited Russia to hack Hillary on nationa"
eprophotog|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: GOP Lobbyist requests AG to investigate Trump for political corruption#cnn #msnbc #AMJoy #cnnsotu #thisweek #res
al_draper|YouTube|0.0|0.0|1.0|0.0|The Rise Of Darth Trump Final: https://t.co/Iz8n37PRF7 via @YouTube
al_draper|youtube|0.0|0.0|1.0|0.0|The Rise Of Darth Trump Final: https://t.co/Iz8n37PRF7 via @YouTube
_flanders|jruha|0.4215|0.0|0.887|0.113|RT @jruha: If this is true #Trump can't be installed. #stribpol #abc #cbs #nbc #cnn #p2 #1u #topprog #Resist #GOP #Fascism #Treason #NoTru
JennHenrichsen|propublica|0.0|0.0|1.0|0.0|How Journalists Need to Go Beyond Fact Checking Trump - ProPublica https://t.co/2qzjDFdWQB via @propublica
JennHenrichsen|propublica|0.0|0.0|1.0|0.0|How Journalists Need to Go Beyond Fact Checking Trump - ProPublica https://t.co/2qzjDFdWQB via @propublica
BettorsChat|MotherJones|0.2023|0.0|0.87|0.13|Donald #Trump  top ten giveaways to Vladimir Putin https://t.co/iy40dDfemx via @MotherJones @BillMaher @MMFlint
BettorsChat|motherjones|0.2023|0.0|0.87|0.13|Donald #Trump  top ten giveaways to Vladimir Putin https://t.co/iy40dDfemx via @MotherJones @BillMaher @MMFlint
SURJColumbusOH|prisonculture|0.2023|0.0|0.904|0.096|RT @prisonculture: Trump's America is just America as it has always existed. I think this is important to know.
Deplorablefrog1|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
POOetryman|Beachfront|-0.6249|0.186|0.814|0.0|RT @Beachfront: @KellyannePolls @ThePressofAC You're a traitor. You're a disaster for your country. You were bought by Trump who is a natio
BemusedDukat|Sargon_of_Akkad|0.34|0.0|0.897|0.103|"@Sargon_of_Akkad The reason Trump speaks bluntly, yet is played 4D chess, is because he's from NY.  That's just how we speak here."
rgrossley48|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
TheKeeper2016|TheDailyEdge|-0.6597|0.253|0.747|0.0|"RT @TheDailyEdge: REMINDER: When asked about Putin killing journalists, Trump equated it w/leadership https://t.co/12C5w9eM8q"
TheKeeper2016|twitter|-0.6597|0.253|0.747|0.0|"RT @TheDailyEdge: REMINDER: When asked about Putin killing journalists, Trump equated it w/leadership https://t.co/12C5w9eM8q"
la__intelectual|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
Bobbyh214|House_Insider|0.5423|0.0|0.774|0.226|RT @House_Insider: https://t.co/Pk8oIA0FD8: We're Going to Start Saying 'Merry Christmas' Again https://t.co/yl8NrxJbyV https://t.co/Vnp2O5
Bobbyh214|twitter|0.5423|0.0|0.774|0.226|RT @House_Insider: https://t.co/Pk8oIA0FD8: We're Going to Start Saying 'Merry Christmas' Again https://t.co/yl8NrxJbyV https://t.co/Vnp2O5
bchek833|HuffPostPol|-0.6192|0.296|0.704|0.0|RT @HuffPostPol: Trump used to complain about Obama not getting intelligence briefings https://t.co/bxEDS3p8yw https://t.co/gWLZe7DoGO
bchek833|m|-0.6192|0.296|0.704|0.0|RT @HuffPostPol: Trump used to complain about Obama not getting intelligence briefings https://t.co/bxEDS3p8yw https://t.co/gWLZe7DoGO
Fooddiva20|TIME|0.0377|0.133|0.727|0.14|"RT @TIME: Donald Trump says he doesn't need daily intelligence briefings because he's a ""smart person"" https://t.co/hE8l3iYAOh"
Fooddiva20|time|0.0377|0.133|0.727|0.14|"RT @TIME: Donald Trump says he doesn't need daily intelligence briefings because he's a ""smart person"" https://t.co/hE8l3iYAOh"
LorenzoQ|ezlusztig|-0.6249|0.17|0.83|0.0|"RT @ezlusztig: Purely on the basis of information publicly available - just the tip of an iceberg, presumably - Obama could devastate Trump"
KatCeccotti|juneday864|0.0|0.0|1.0|0.0|"RT @juneday864: Um, I am 100% concerned Trump, and everyone propping him up, is an unapologetic traitor. https://t.co/DGhCSQZBaL"
KatCeccotti|twitter|0.0|0.0|1.0|0.0|"RT @juneday864: Um, I am 100% concerned Trump, and everyone propping him up, is an unapologetic traitor. https://t.co/DGhCSQZBaL"
ProAssad|ABC|0.2023|0.197|0.574|0.23|"RT @ABC: Where Trump's critics see conflicts of interest, his global business partners see opportunities. @brianross reports: https://t.co/"
ProAssad|t|0.2023|0.197|0.574|0.23|"RT @ABC: Where Trump's critics see conflicts of interest, his global business partners see opportunities. @brianross reports: https://t.co/"
JHSaunders|AP|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
JHSaunders|t|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
BlameThe1st|Nash076|-0.5574|0.122|0.878|0.0|"RT @Nash076: By all means, explain to your 10 year old that they don't get to see Star Wars because the writers were mean to Trump. #DumpSt"
browntom1234|dem_happy|-0.4926|0.259|0.741|0.0|@dem_happy It's what Satan uses to dupe cucks into disobeying or questioning emperor Trump!
lolife52|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
lolife52|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
CDCollector23|gunsrus7|0.0|0.0|1.0|0.0|@gunsrus7 Trump is nothing more than an overgrown Putin puppet because he owes his entire election to Russian interference.
PiratesWife82|Will_Bunch|-0.7149|0.239|0.761|0.0|"RT @Will_Bunch: Worse than Watergate? Russia hacking is massive cloud over Trump presidency, and America. What caused this big mess? https:"
Kim38875219|CNBC|0.0|0.0|1.0|0.0|"RT @CNBC: Trump says U.S. not necessarily bound by ""one China"" policy https://t.co/hkRFMZLkxO"
Kim38875219|cnbc|0.0|0.0|1.0|0.0|"RT @CNBC: Trump says U.S. not necessarily bound by ""one China"" policy https://t.co/hkRFMZLkxO"
CaroleMyers|McJesse|0.0|0.0|1.0|0.0|RT @McJesse: We thought Trump was Tweeting in middle of the night. Now we know he's just on Moscow time.
Jude5253|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
anicho47|LibAmericaOrg|-0.3254|0.127|0.873|0.0|RT @LibAmericaOrg: SHOCKER: Russias Head Of Foreign Affairs Thinks Trumps Sec Of State Pick Is Awesome(Tweets) https://t.co/ETCe0GYtPk
anicho47|liberalamerica|-0.3254|0.127|0.873|0.0|RT @LibAmericaOrg: SHOCKER: Russias Head Of Foreign Affairs Thinks Trumps Sec Of State Pick Is Awesome(Tweets) https://t.co/ETCe0GYtPk
PubPolHist|DLin71|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
PubPolHist|twitter|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
Ximeko|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
MiaEvan30311368|johndurant|-0.25|0.233|0.6|0.167|RT @johndurant: Wealthy Hollywood celebrity assaults Uber driver over Trump: https://t.co/nM4eXaGKLa
MiaEvan30311368|deadline|-0.25|0.233|0.6|0.167|RT @johndurant: Wealthy Hollywood celebrity assaults Uber driver over Trump: https://t.co/nM4eXaGKLa
debyoungblood|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
breakfastqueen1|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
modernbob|WSJ|0.0772|0.12|0.705|0.174|"RT @WSJ: Defending his recent attacks on corporate America, Trump said: I want us to make good deals for this countryhttps://t.co/yUgF9S"
DickNixonLives|Evan_McMullin|0.0|0.0|1.0|0.0|@Evan_McMullin @realDonaldTrump face it Evan you have been begging Trump for a cabinet post the whole time
LindaWestbroo11|NormEisen|0.595|0.101|0.668|0.231|"RT @NormEisen: Wow, Trump has just 41% approval (vs 72 at this pt 4 Obama) with 65% concerned that his business ties CONFLICT. https://t.co"
LindaWestbroo11|t|0.595|0.101|0.668|0.231|"RT @NormEisen: Wow, Trump has just 41% approval (vs 72 at this pt 4 Obama) with 65% concerned that his business ties CONFLICT. https://t.co"
studygoddess01|law_newz|-0.5267|0.236|0.764|0.0|Melania Trump's 'Revenge Lawyer' Apparently Doesn't Understand First Amendment https://t.co/RJ2tCKaWXc via @law_newz
studygoddess01|lawnewz|-0.5267|0.236|0.764|0.0|Melania Trump's 'Revenge Lawyer' Apparently Doesn't Understand First Amendment https://t.co/RJ2tCKaWXc via @law_newz
NewsdeskUS|bbc|0.0|0.0|1.0|0.0|Trump on Twitter https://t.co/XqxeeDIEIm
TheMrsDarcy|laurie6805|0.0|0.0|1.0|0.0|RT @laurie6805: https://t.co/meA70vnfVt
TheMrsDarcy|dailycaller|0.0|0.0|1.0|0.0|RT @laurie6805: https://t.co/meA70vnfVt
messerduff|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
ChristineAdams3|DataLogicTruth|0.6305|0.101|0.594|0.305|"RT @DataLogicTruth: Trump says he doesn't need intelligence briefings because ""I'm, like, a smart person.""We can all agree: false premise"
lovemedietcoke|tonyschwartz|-0.296|0.091|0.909|0.0|RT @tonyschwartz: I don't believe anything Donald Trump says. Not one word. It is all manipulation and mind games all the time. (Same for K
DessyFenix|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: Now - with Trump as the non-conformist, not-like-all-the-other-rotten-conspiratorial-assholes paragon, the Russians go int"
inklake|France4Hillary|-0.4514|0.217|0.616|0.167|RT @France4Hillary: It makes me SO SICK to see that Trump is lying about the Russian help he received to win the election. MAN UP &amp; TELL TH
breaguiniga|Laughbook|0.0|0.0|1.0|0.0|RT @Laughbook: Even Barron Trump don't believe in his dad Donald Trump https://t.co/yK5Rp8EDH1
breaguiniga|twitter|0.0|0.0|1.0|0.0|RT @Laughbook: Even Barron Trump don't believe in his dad Donald Trump https://t.co/yK5Rp8EDH1
kaleemarie24|feliciaw5853|-0.2263|0.148|0.742|0.109|"RT @feliciaw5853: Obama trapped in presidency defining moment. Like Lincoln, unavoidable decision. Have CIA release intel on Trump. https:/"
kaleemarie24||-0.2263|0.148|0.742|0.109|"RT @feliciaw5853: Obama trapped in presidency defining moment. Like Lincoln, unavoidable decision. Have CIA release intel on Trump. https:/"
KathyFeingold|TheDailyEdge|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
KathyFeingold|twitter|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
EdouardDugas|Claude2052|0.0|0.0|1.0|0.0|Time to go back to school.@Claude2052 #polqc #polcan #rnc #gop #trump https://t.co/vxsNcRZlLc
EdouardDugas|twitter|0.0|0.0|1.0|0.0|Time to go back to school.@Claude2052 #polqc #polcan #rnc #gop #trump https://t.co/vxsNcRZlLc
MythicalStig|markmobility|-0.3612|0.135|0.865|0.0|RT @markmobility: NYT Editorial: On Trump's refusal to investigate Russia. The election was indeed rigged. https://t.co/aRKMthkimV https://
MythicalStig|nytimes|-0.3612|0.135|0.865|0.0|RT @markmobility: NYT Editorial: On Trump's refusal to investigate Russia. The election was indeed rigged. https://t.co/aRKMthkimV https://
trudgintheroad|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
Stephan19330818|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
PattiPropst|breitbart|0.0|0.0|1.0|0.0|https://t.co/xzTse7iztU
KathyTu57558497|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
KathyTu57558497|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
DonMcKenzie|Delo_Taylor|-0.3818|0.094|0.906|0.0|"RT @Delo_Taylor: If the goal was to keep Trump from ever becoming POTUS, the first thing you shoulda done was fight to keep HRC from being"
vandives|mtracey|-0.5423|0.268|0.632|0.1|"RT @mtracey: Yes, stake your opposition to Trump on CIA hearsay, treason accusations, and Russia paranoia. More sound strategic thinking fr"
hypnocoach183|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
hypnocoach183|change|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
TerryGomez91|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
DRHsPsychoCafe|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
Lina_J_Al|Joyce_Karam|-0.8176|0.309|0.691|0.0|RT @Joyce_Karam: There's an attack on Church in Egypt;Terror in Istanbul; ISIS took Palmyra; CIA alarm on Russia.But #Trump is attacking NB
andersongouldjr|DeanLeh|0.4939|0.0|0.862|0.138|RT @DeanLeh: 5 million Americans sign the petition to the Electoral College begging them to save us from the Trump NIGHTMARE: https://t.co/
andersongouldjr|t|0.4939|0.0|0.862|0.138|RT @DeanLeh: 5 million Americans sign the petition to the Electoral College begging them to save us from the Trump NIGHTMARE: https://t.co/
DKWilson56|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
faabbbs|BraddJaffy|-0.5994|0.218|0.782|0.0|RT @BraddJaffy: President Obama and President-elect Trump react to the death of Fidel Castro https://t.co/Teg8dA4D7e
faabbbs|twitter|-0.5994|0.218|0.782|0.0|RT @BraddJaffy: President Obama and President-elect Trump react to the death of Fidel Castro https://t.co/Teg8dA4D7e
AnnaHarffey|DataLogicTruth|0.4588|0.094|0.684|0.222|"RT @DataLogicTruth: Trump: ""From everything I see, Putin has no respect for this person.""Clinton: ""Well thats because he'd rather have a"
neighborlee|DeAnnSmithkc|0.0|0.0|1.0|0.0|@DeAnnSmithkc @SallyAlbright Comey &amp; rallies where trump attempts #incite2riot my fingernail has more class/morals .
RayREllis1|YouTube|0.0|0.0|1.0|0.0|"Trump ""AMERICA"": https://t.co/66MP9QeyCA via @YouTube"
RayREllis1|youtube|0.0|0.0|1.0|0.0|"Trump ""AMERICA"": https://t.co/66MP9QeyCA via @YouTube"
sp1ritharambe|ananavarro|0.0|0.0|1.0|0.0|@ananavarro Ana had to get that one Trump dig in.. Part of her contract at CNN.
ccbean1965|steph93065|-0.4019|0.112|0.843|0.044|"RT @steph93065: Until Jan 20, the left/MSM will do/say anything to delegitimize &amp; try to prevent Trump from taking office; their tantrum is"
lolalolita0|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/TEGHqhLpZN https://t.co"
lolalolita0|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/TEGHqhLpZN https://t.co"
VictorMoruzzi|BBCWorld|0.0|0.0|1.0|0.0|RT @BBCWorld: Trump on Twitter https://t.co/RCADyEifSU
VictorMoruzzi|bbc|0.0|0.0|1.0|0.0|RT @BBCWorld: Trump on Twitter https://t.co/RCADyEifSU
79topper|JoyAnnReid|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
79topper|twitter|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
val_kudirka|cleo_peterson|-0.6027|0.304|0.696|0.0|RT @cleo_peterson: #TrumpIsTreason #NotMyPresident #NotMyCountry Charge Trump with TREASON! https://t.co/Ozqzr6wmRk
val_kudirka|twitter|-0.6027|0.304|0.696|0.0|RT @cleo_peterson: #TrumpIsTreason #NotMyPresident #NotMyCountry Charge Trump with TREASON! https://t.co/Ozqzr6wmRk
nigelcameron|20committee|0.2023|0.0|0.924|0.076|RT @20committee: Trump's refusal to admit that Russia was behind election games is forcing his cabinet nominees to lie publicly in ways the
93skedoo|Fusion|0.0|0.0|1.0|0.0|@Fusion but it's not news it's propoganda and it's been a concerted campaign https://t.co/rFHFsl20eY
93skedoo|theguardian|0.0|0.0|1.0|0.0|@Fusion but it's not news it's propoganda and it's been a concerted campaign https://t.co/rFHFsl20eY
LaOkieKat|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
LaOkieKat|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
It_is_NunyaDB|Fusion|-0.7003|0.279|0.721|0.0|RT @Fusion: This CNN segment shows just how big of a problem fake news has become: https://t.co/fvPIgcGtJu https://t.co/FLo8C3k7iv
It_is_NunyaDB|fusion|-0.7003|0.279|0.721|0.0|RT @Fusion: This CNN segment shows just how big of a problem fake news has become: https://t.co/fvPIgcGtJu https://t.co/FLo8C3k7iv
allthatyaaazzzz|business|0.0|0.0|1.0|0.0|RT @business: Trump's businesses made more than $14.6 million off of his campaign https://t.co/YDwtF3KW8Z https://t.co/7NWdmyaoUV
allthatyaaazzzz|bloomberg|0.0|0.0|1.0|0.0|RT @business: Trump's businesses made more than $14.6 million off of his campaign https://t.co/YDwtF3KW8Z https://t.co/7NWdmyaoUV
lindsayrda53|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/Z7ruXdiBFu https://t.co/j1GAYDRau5
lindsayrda53|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/Z7ruXdiBFu https://t.co/j1GAYDRau5
Rajivkapoor2318|Newsmax|-0.7003|0.326|0.674|0.0|Michael Moore Plans to Protest at Trump Inauguration https://t.co/NLYMXzYmVq via @Newsmax moore looks obscene
Rajivkapoor2318|newsmax|-0.7003|0.326|0.674|0.0|Michael Moore Plans to Protest at Trump Inauguration https://t.co/NLYMXzYmVq via @Newsmax moore looks obscene
DanielMichaelJ|DLin71|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
DanielMichaelJ|twitter|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
McbrideHoover|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
ArtHauntsMe|EJR91372|-0.2023|0.131|0.766|0.102|@EJR91372 lol. It's not that covert. It just means everyone is digging up old shit about Trump's visits and dealing with the Russkies
diannabythesea|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
l8j42|cia|-0.0772|0.134|0.746|0.119|.@cia @FBI i will gladly hear the secrets trump is refusing to hear LMK where to sign up
Markus03121966|BrendanNyhan|0.0|0.0|1.0|0.0|"RT @BrendanNyhan: Trump: ""I am turning down billions of dollars of deals."" Oh?"
PamelafBrockman|mateagold|-0.296|0.121|0.879|0.0|RT @mateagold: No president in recent history has filled a Cabinet with so many major donors. https://t.co/BbnJC608JZ https://t.co/zX9UKLSL
PamelafBrockman|washingtonpost|-0.296|0.121|0.879|0.0|RT @mateagold: No president in recent history has filled a Cabinet with so many major donors. https://t.co/BbnJC608JZ https://t.co/zX9UKLSL
ChoocfantasyM|tonyschwartz|-0.296|0.091|0.909|0.0|RT @tonyschwartz: I don't believe anything Donald Trump says. Not one word. It is all manipulation and mind games all the time. (Same for K
scutify|scutify|0.0|0.0|1.0|0.0|Bi-Weekly Economic Review: Trump Catches A Tailwind https://t.co/CWcZ8gqvte $USD $GOLD $IWM #bonds #commodities #credit #spreads #dollar
IntrovertRN1975|JuddLegum|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
IntrovertRN1975|medium|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
undercover0000|shareblue|-0.5499|0.258|0.621|0.12|Kellyanne Conway says Trump is going to put his own people in the intelligence community https://t.co/0gpaHFJLsy      NUTS! Just NUTS!
catlover1943|CDZ_999|-0.8828|0.339|0.661|0.0|RT @CDZ_999: i just heard trump say he doesnt want to sit thru them . get this fuck outta contention or you are DOOMED https://t.co/3Xgk0HF
catlover1943|t|-0.8828|0.339|0.661|0.0|RT @CDZ_999: i just heard trump say he doesnt want to sit thru them . get this fuck outta contention or you are DOOMED https://t.co/3Xgk0HF
Presley48R|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
Presley48R|thegatewaypundit|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
bethtomkiw|mradamscott|0.7345|0.0|0.721|0.279|"RT @mradamscott: In short our president-elect, in cahoots with Russia, seems determined on dismantling our republic. Merry Christmas!https"
Michell66010778|amjoyshow|0.0|0.0|1.0|0.0|RT @amjoyshow: .@JoyAnnReid just explained all the people linked to Donald Trump who have documented ties to #Russia and Putin #AMJoy https
YoyoStube|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
elisabetta7991|YourAnonCentral|0.0|0.0|1.0|0.0|RT @YourAnonCentral: Democracy doesn't trump human rights. @DrHaque
APOYODECHILE|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
RegaloDelSenor|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
zumausa|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
HondaMashburn|CapehartJ|0.0|0.0|1.0|0.0|"RT @CapehartJ: In less than 5 weeks, Trump has revealed just how fragile the Constitution is. https://t.co/DG9Yiz5SYL"
HondaMashburn|washingtonpost|0.0|0.0|1.0|0.0|"RT @CapehartJ: In less than 5 weeks, Trump has revealed just how fragile the Constitution is. https://t.co/DG9Yiz5SYL"
nancy73gg|andieiamwhoiam|0.5267|0.065|0.75|0.185|"RT @andieiamwhoiam: Sorry Lefties, Russians, recounts, aliens (the extraterrestrial kind)...you will never get a new election.  Trump won."
Myocz|Lettradus|-0.296|0.167|0.833|0.0|"RT @Lettradus: ""No sou Politicamente Correto, prefiro ser Honesto"" - Donald Trump https://t.co/MsGWiOSGBn"
Myocz|twitter|-0.296|0.167|0.833|0.0|"RT @Lettradus: ""No sou Politicamente Correto, prefiro ser Honesto"" - Donald Trump https://t.co/MsGWiOSGBn"
PatPatojson|Zeke311|-0.5707|0.185|0.749|0.066|RT @Zeke311: 'The Trump Way': Exclusive Interview Break Down  Alex Jones' Infowars: There's a war on for your mind! https://t.co/lWTGkdpYbY
PatPatojson|infowars|-0.5707|0.185|0.749|0.066|RT @Zeke311: 'The Trump Way': Exclusive Interview Break Down  Alex Jones' Infowars: There's a war on for your mind! https://t.co/lWTGkdpYbY
cvasilevski|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
cvasilevski|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
johnnymercerfan|DLin71|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
johnnymercerfan|twitter|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
carpet_bomber|WSJ|0.0772|0.12|0.705|0.174|"RT @WSJ: Defending his recent attacks on corporate America, Trump said: I want us to make good deals for this countryhttps://t.co/yUgF9S"
maluza56|QuadratinMexico|0.0|0.0|1.0|0.0|"RT @QuadratinMexico: Ante incertidumbre por Trump, hay que promover consumo local: Glvez  https://t.co/4FEiOYmyYR"
maluza56|mexico|0.0|0.0|1.0|0.0|"RT @QuadratinMexico: Ante incertidumbre por Trump, hay que promover consumo local: Glvez  https://t.co/4FEiOYmyYR"
debyoungblood|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
djgirl40|AlecBaldwin|0.9208|0.0|0.516|0.484|"So @AlecBaldwin won for best guest appearance for @nbcsnl...guess his Trump impression wasn't so bad afterall, huh @realDonaldTrump.#SNL"
tobyonekonobe|surfermom77|-0.4215|0.128|0.872|0.0|"RT @surfermom77: The GOP bitter traitors &amp; Estab hacks, McCain &amp; Graham are joining Dems pushing the hairbrained #RussianHacking plothttps"
efox17|FrankLuntz|0.5261|0.0|0.82|0.18|"RT @FrankLuntz: Sometimes, the facts will be favorable to Trump Sometimes, they won't be.But don't only pay attention to the facts that"
andrea_manea|davidfrum|0.7351|0.0|0.754|0.246|"RT @davidfrum: US intelligence community: Russia acted to install Trump. 18 months from now, there wont be a US intelligence community wor"
nice2bcalm|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
nice2bcalm||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
plowman_robert|mikandynothem|0.3802|0.088|0.767|0.146|RT @mikandynothem: Ruth Bader Ginsburg said she would resign if Trump won. Hit the road lady! That will give Trump even more Conservatives
Lewisgd|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
Damuhar|lulach_cuardach|0.0|0.0|1.0|0.0|RT @lulach_cuardach: @Slender_Sir @nydwracu That little boy's name?Donald J. Trump.
whaaf|Adenovir|-0.8658|0.386|0.614|0.0|"RT @Adenovir: Carl Bernstein, who broke the Watergate scandal that led to Nixon's resignation, said that Nixon's lies were nothing compared"
dashing_reaver|_premiumfan|-0.6124|0.192|0.808|0.0|@_premiumfan @BillNemacheck It sucks when you find out how much Trump sucks and how he's MORE corrupt and you still voted for him
respectinc|jayrosen_nyu|0.4168|0.0|0.878|0.122|"RT @jayrosen_nyu: 3/ There, the implied message from journalism to the Trump forces (the government + his core supporters) is: ""Don't hurt"
TWalterErickson|JoeBerkowitz|0.0|0.0|1.0|0.0|RT @JoeBerkowitz: This is the most patriotic thing an American can do right now. https://t.co/htXS14yRlA
TWalterErickson|politico|0.0|0.0|1.0|0.0|RT @JoeBerkowitz: This is the most patriotic thing an American can do right now. https://t.co/htXS14yRlA
ltwhite|thehill|0.0|0.0|1.0|0.0|RT @thehill: Trump goes after NBC news in tweethttps://t.co/32I8myfDsw https://t.co/vj13vixfUJ
ltwhite|twitter|0.0|0.0|1.0|0.0|RT @thehill: Trump goes after NBC news in tweethttps://t.co/32I8myfDsw https://t.co/vj13vixfUJ
joh53293471|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
usmaan_aisha|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
jzd3|nbcsnl|0.0|0.0|1.0|0.0|RT @nbcsnl: BREAKING: President-elect Trump picks Walter White as Head of DEA. https://t.co/h3EtN3QFQO #CenaOnSNL https://t.co/vuJPKIsYqM
jzd3|nbc|0.0|0.0|1.0|0.0|RT @nbcsnl: BREAKING: President-elect Trump picks Walter White as Head of DEA. https://t.co/h3EtN3QFQO #CenaOnSNL https://t.co/vuJPKIsYqM
Adriene26|yashar|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
Adriene26|twitter|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
grandpooba5440|rudepundit|-0.5719|0.207|0.712|0.081|RT @rudepundit: Trump made the Russia story worse by attacking the CIA. An innocent man would have stated his concern and called for invest
SRStalcup|thehill|-0.6305|0.232|0.768|0.0|"@thehill post hoc, ergo propter hoc. The country is stuck with Trump and Clinton wasn't that super anyroad. Lose/lose."
INSOMNIAK_DJ|HamiltonElector|0.2298|0.123|0.757|0.12|"RT @HamiltonElector: Mr. Trump you are hardly a genius, no matter what Comrade Putin says.  We are smarter than you. We are #hamiltonelecto"
jen_thorson|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
Inked1BNA|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
Inked1BNA|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
lsuagain|PSheritaakkloh|-0.6199|0.238|0.762|0.0|"@PSheritaakkloh @manuufs If you hate Trump, why are you following his tweets? Troll much?"
Chi_Ship|soit_goes|0.8225|0.0|0.752|0.248|.@soit_goes does the trump win equate to the Mittens win in 2012? Will the @realDonaldTrump take the US to its knees and start the uprising.
tonic516|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Ltr from Hon Elijah Cummings asking Chaffetz to Investigate Trump biz conflicts#cnn #msnbc #AMJoy #cnnsotu #this
AtlTeaPartyLove|twitter|-0.0572|0.071|0.929|0.0|Women that voted for Trump used their brain.They didn't want a president just because she has a vagina. https://t.co/MQdEUpvOJN
anthonygbrooks|twitter|0.4404|0.0|0.873|0.127|"If 500 Trump supporters rally in Boston I'll cover them, 2. Btw, u shd learn the diff between PBS &amp; NPR https://t.co/0szbd1sf51"
IntrovertRN1975|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 7. Therefore, it could be a ""false flag"" operation by the Obama administration https://t.co/oRUPSkz7NV"
IntrovertRN1975|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 7. Therefore, it could be a ""false flag"" operation by the Obama administration https://t.co/oRUPSkz7NV"
JenTromans|CaptainsLog2016|-0.0258|0.064|0.936|0.0|RT @CaptainsLog2016: Funneling millions in campaign $ to his businessesSelling Cabinet positions &amp; MAGA hatsTrump may actually become a
Kashinka|Endoraknows|0.4891|0.118|0.673|0.209|RT @Endoraknows: @wvjoe911 I agree !! Why pay ours when Trump doesn't pay his? No taxation without representation- Trump doesn't represent
Bayathread|HuffPostWomen|0.5859|0.0|0.703|0.297|@HuffPostWomen follow @RachelleHodgs for brilliant graphing of Trump word salads.
julstitt|realDonaldTrump|0.636|0.102|0.625|0.273|"@realDonaldTrump Trump has jumped in the swamp to take from the poor. Research his cabinet staff, only out to benefit wealthy, like himself!"
brianpiero|Deanofcomedy|-0.2732|0.1|0.9|0.0|RT @Deanofcomedy: .@petemont of @peoplefor talks on my  @SXMInsight show about risk of Christian Dominionism in America under Trump: https:
Shanny_resqchi|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
trungngo09|georgebkk|0.0772|0.0|0.86|0.14|RT @georgebkk: Thailand awaits Trumps foreign policy team https://t.co/teJ5BMrLNh
trungngo09|thaivisa|0.0772|0.0|0.86|0.14|RT @georgebkk: Thailand awaits Trumps foreign policy team https://t.co/teJ5BMrLNh
washumom|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: New York Times Editorial Board demands Donald Trump go along with Russia investigation https://t.co/Fv74uavXcI via @dailynew
washumom|dailynewsbin|0.0|0.0|1.0|0.0|RT @starfirst: New York Times Editorial Board demands Donald Trump go along with Russia investigation https://t.co/Fv74uavXcI via @dailynew
thebobbyb|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
notastalker_uR|nbcsnl|0.4588|0.0|0.769|0.231|"RT @nbcsnl: Welcome to the Trump administration, Walter White. #CenaOnSNL https://t.co/aPaceUQcO0"
notastalker_uR|twitter|0.4588|0.0|0.769|0.231|"RT @nbcsnl: Welcome to the Trump administration, Walter White. #CenaOnSNL https://t.co/aPaceUQcO0"
eprophotog|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Ltr from Hon Elijah Cummings asking Chaffetz to Investigate Trump biz conflicts#cnn #msnbc #AMJoy #cnnsotu #this
xfigmentx|Khanoisseur|-0.4588|0.15|0.85|0.0|RT @Khanoisseur: 2 reasons for trump rejecting daily intel briefings:1. Plausible deniability2. Busy making side deal$$ for himself @mrp
nettsarie|TeenVogue|0.0|0.0|1.0|0.0|Donald Trump Is Gaslighting America https://t.co/RFqtn75HnJ via @TeenVogue
nettsarie|teenvogue|0.0|0.0|1.0|0.0|Donald Trump Is Gaslighting America https://t.co/RFqtn75HnJ via @TeenVogue
jennifer4nm|kurteichenwald|-0.5423|0.176|0.824|0.0|"RT @kurteichenwald: Fox/Cheney went nuts when found out Obama got intel briefings in writing, rather than read to him. But Trump no briefin"
cdat|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Hellon_Heels|SpeakerRyan|-0.296|0.109|0.891|0.0|.@SpeakerRyan Trump &amp; his Russia ties are a #StateofEmergency. Sign a letter from the people to stop Trump Jan. 6. https://t.co/raNLdFh810
Hellon_Heels|npr|-0.296|0.109|0.891|0.0|.@SpeakerRyan Trump &amp; his Russia ties are a #StateofEmergency. Sign a letter from the people to stop Trump Jan. 6. https://t.co/raNLdFh810
ZiggyinHeavon|redstatewatcher|-0.5983|0.393|0.607|0.0|Boom! Trump destroys NBC Nightly News https://t.co/0Com4mGiTY
demfemme|pittgriffin|0.2654|0.117|0.674|0.21|RT @pittgriffin: Trump's poodles don't care.'Chris Wallace Confronts #Trump on Conflicts of Interest: You Hammered Hillary Clinton' https
KHZ4HGP|aol|-0.3311|0.469|0.192|0.339|LOL! Oh Hell. https://t.co/zlVJaxihec
shhendrickson|surfermom77|-0.4215|0.128|0.872|0.0|"RT @surfermom77: The GOP bitter traitors &amp; Estab hacks, McCain &amp; Graham are joining Dems pushing the hairbrained #RussianHacking plothttps"
PizzaAbuser|sherlockmichael|-0.296|0.25|0.593|0.157|RT @sherlockmichael: Trump voters:Has confirmation of Russia's illegal role in Trump's success made you skeptical of a #TrumpPresidency?
wikkidwillow|SenSanders|0.2023|0.058|0.853|0.089|RT @SenSanders: Mr. Trump told working people he was on their side. Millions of us are going to demand that he keep his promise.
sampson_elaine|DailyNewsBin|0.4767|0.0|0.829|0.171|RT @DailyNewsBin: Intelligence community fires back at Donald Trump after he dismisses CIAs Russia findings https://t.co/LsmDQAulB6
sampson_elaine|dailynewsbin|0.4767|0.0|0.829|0.171|RT @DailyNewsBin: Intelligence community fires back at Donald Trump after he dismisses CIAs Russia findings https://t.co/LsmDQAulB6
Luvnstuff2|thr|0.0|0.0|1.0|0.0|Michael Moore Details Plans for Trump's Inauguration https://t.co/F0tHNWka8p via @thr
Luvnstuff2|hollywoodreporter|0.0|0.0|1.0|0.0|Michael Moore Details Plans for Trump's Inauguration https://t.co/F0tHNWka8p via @thr
ProAssad|nytimesworld|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
ProAssad|nytimes|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
danni_rie|JuddLegum|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
danni_rie|t|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
AmazingAshesly|elijahdaniel|0.8109|0.0|0.731|0.269|RT @elijahdaniel: MY FRIEND WAS AT THE WHITE HOUSE CHRISTMAS PARTY AND ASKED FUCKING BARACK OBAMA WHAT HE THOUGHT ABOUT TRUMP TEMPTATIONS I
euphoricpieta|TheThomason|0.0|0.0|1.0|0.0|"RT @TheThomason: Realistically, I just don't know if there's time for Trump to learn to read before beginning his presidency."
suicide_romance|Hellon_Heels|0.0|0.0|1.0|0.0|RT @Hellon_Heels: #Leninist Trump and Bannon r traitors #StopTrump https://t.co/5tZArlpOP3
suicide_romance|twitter|0.0|0.0|1.0|0.0|RT @Hellon_Heels: #Leninist Trump and Bannon r traitors #StopTrump https://t.co/5tZArlpOP3
SturdeeBeggar|_0HOUR1|-0.5574|0.187|0.813|0.0|RT @_0HOUR1: Trump should also cut all of John McCain foreign fighting money immediately @realDonaldTrump That is what its about the billio
Jeff_Leader|ericgarland|-0.529|0.189|0.811|0.0|RT @ericgarland: The Russians didn't create Trump - only New York City and American gullibility could have done that.But they've got a SW
breakfastqueen1|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
ArianeBellamar|TheJusticeDept|0.0|0.0|1.0|0.0|#ARRESTTRUMP Calling on the @TheJusticeDept to #prosecute #Trump! #RESIST #RussiaHacking #sexism #racism #LockHimUp https://t.co/D1U76dohrZ
ArianeBellamar|change|0.0|0.0|1.0|0.0|#ARRESTTRUMP Calling on the @TheJusticeDept to #prosecute #Trump! #RESIST #RussiaHacking #sexism #racism #LockHimUp https://t.co/D1U76dohrZ
websterwakeemup|SocialPowerOne1|-0.0772|0.254|0.565|0.181|@SocialPowerOne1 There will be many peaceful protests because Trump has lied so often.
Tuscan21_PM|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
soaksponge|MichaelDelauzon|0.0|0.0|1.0|0.0|RT @MichaelDelauzon: Secret Service nabs Ivanka Trump's stalker for the second time. Justin Massler busted last May and again this week. ht
MtLion15|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
MtLion15||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
ShutUpBabyINoIt|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
RichardTrubacek|thehill|0.0|0.0|1.0|0.0|Trump lashes out at NBC News on Twitter https://t.co/y63SjN08iK
EnriqueM77|WG_Burton|0.1531|0.0|0.833|0.167|RT @WG_Burton: A Carefully Planned Operation to Prevent President-elect Donald Trumps Accession to the White House?https://t.co/HQHpFUBoH
EnriqueM77|t|0.1531|0.0|0.833|0.167|RT @WG_Burton: A Carefully Planned Operation to Prevent President-elect Donald Trumps Accession to the White House?https://t.co/HQHpFUBoH
KangJiaChen|tomphillipsin|-0.7783|0.264|0.736|0.0|"RT @tomphillipsin: Beijing life, late 2016: wake up, inhale smog, think, 'What the hell did Donald Trump say while I was sleeping?'"
ValkyrieSigrid|US_Army_Vet|0.3716|0.0|0.846|0.154|RT @US_Army_Vet: Judge Napolitano: NSA not Russia hacked Hillary! Judge Jeanine Slams Obamahttps://t.co/Tzykej89gp @LeahR77 #USAhttps:
winkiechance|Bane1349|-0.128|0.145|0.727|0.127|RT @Bane1349: Indeed.. We would follow President Trump To Hell... And BackZero Loyalty to Them.  Just look at those two Bastards Graham M
waldmania|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
tedreally|yashar|0.6808|0.0|0.772|0.228|@yashar And yet none of them use language that attracts Trump supporters. When will they learn to use his language style?
peggyhsinhsin|TeenVogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
peggyhsinhsin|teenvogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
ramrhonda|sjredmond|-0.7269|0.253|0.747|0.0|RT @sjredmond: I don't think Trump will ever get to #MAGA. His schtick is all #MARS: Make America Rude &amp; Selfish.
amerycarlson|WayneDupreeShow|-0.4767|0.171|0.829|0.0|RT @WayneDupreeShow: Rep. Tulsi Gabbard Says Democrats Wrong To Bash Trump For Retired General Picks https://t.co/62oDMIBBmO
amerycarlson|newsninja2012|-0.4767|0.171|0.829|0.0|RT @WayneDupreeShow: Rep. Tulsi Gabbard Says Democrats Wrong To Bash Trump For Retired General Picks https://t.co/62oDMIBBmO
SammyMorgan91|nytimes|0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
SammyMorgan91||0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
EllyHuy|youtube|-0.5574|0.223|0.777|0.0|Ti  thm video vo danh sch pht https://t.co/LjhP6mX323 WIKILEAKS FBI NEWS: Trumps FBI Probe Contradicts CIA. No Link
texlaker|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
as_promised|addictinginfo|-0.1027|0.142|0.733|0.125|Are Trump Supporters Too Dumb To Know Theyre Dumb?Science Says Probably https://t.co/GxytTqA0Xv &lt;or to know what #DunningKruger effect is
PIE20121|yashar|-0.4215|0.149|0.851|0.0|@yashar @StillLes4Hill And yet Carl Bernstein enabled Trump to happen with his lies and smears of HRC.
jtmcfluffy|DLin71|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
jtmcfluffy|twitter|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
BVenditte|AriMelber|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
BVenditte|t|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
JohnSede|NewsBud_|0.0|0.0|1.0|0.0|RT @NewsBud_: #Trump Fills the Swamp With Steven Mnuchin https://t.co/GQHmeCjT4h https://t.co/B5NNaN2NIF
JohnSede|boilingfrogspost|0.0|0.0|1.0|0.0|RT @NewsBud_: #Trump Fills the Swamp With Steven Mnuchin https://t.co/GQHmeCjT4h https://t.co/B5NNaN2NIF
KathyLangeNovak|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
Tenkellers|RedNationRising|-0.6808|0.235|0.765|0.0|RT @RedNationRising: HIDDEN CAM: Professor Says Trump Election an 'Act of Terrorism' #RedNationRising  https://t.co/BJDNT0FQSD via @scrowder
Tenkellers|louderwithcrowder|-0.6808|0.235|0.765|0.0|RT @RedNationRising: HIDDEN CAM: Professor Says Trump Election an 'Act of Terrorism' #RedNationRising  https://t.co/BJDNT0FQSD via @scrowder
777Francejacque|V_of_Europe|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
777Francejacque|thegatewaypundit|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
journeysincolor|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
Camilian1Sabel|RichardTBurnett|0.8316|0.0|0.63|0.37|RT @RichardTBurnett: Everything is coming back thanks to Donald Trump:1. Pride in America.2. Saluting American flag.3. Merry Christmas.
Mandari25733571|girlsreallyrule|0.4648|0.0|0.888|0.112|"RT @girlsreallyrule: The CIA is SURE Russia helped elect Trump, the FBI is not as sure...Hmmm. One of these things is Comey-er than the oth"
sarge19k4088|CarlaChamorros|0.0|0.0|1.0|0.0|"RT @CarlaChamorros: Vintage Trump, listen and understand why HE/WE WON:Exclusive: Donald Trump on Cabinet picks, transition process https"
AlekseiTheWolf|marling981|0.7096|0.084|0.602|0.314|@marling981 @CoryBooker Seems like a good idea til you realize that people will want to clean up the mess left after Trump's bubble pops
leilacountry|yolandazavala7|-0.296|0.167|0.833|0.0|@yolandazavala7 fbi report says no russian associated with trump or his associates
MaryTrinetti|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
_missnher|twitter|0.0|0.0|1.0|0.0|Trump https://t.co/GiTfFNY2sA
DtRh321|Yvette_G_Nacer|0.4588|0.0|0.571|0.429|"@Yvette_G_Nacer trump's ""russian"" server. haha"
ABSFSU1|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
respectinc|jayrosen_nyu|0.2732|0.0|0.913|0.087|RT @jayrosen_nyu: 2/ Already in gear: Trump loyalists (Jeffrey Lord is the model) recruited into the press as a gaudy show of balance. http
TechNewsDB|technewsdb|0.0|0.0|1.0|0.0|"Larry Page, Tim Cook said to attend Donald Trump's tech summit     - CNET - https://t.co/qf48qX58P4 https://t.co/2DXQBT8h3G"
dblair54|carlreiner|-0.34|0.208|0.66|0.132|"RT @carlreiner: As elated as I was about seeing Dick Van Dyke Show In color tonite, that's how depressed I am about Trump's choices for U.S"
politicsrecycle|teaparty|-0.7154|0.374|0.626|0.0|EXPOSED  Look Whos Behind Scheme to STEAL Trumps Electoral College Votes   https://t.co/3mVyOnVwMu
michaeldhensel|gizmodo|0.0|0.0|1.0|0.0|Finally a plan from Trump. https://t.co/IuvJhJ8HdT
Newyorker2212|DerronDjjrdn|-0.4939|0.167|0.833|0.0|RT @DerronDjjrdn: Donald Trump Keeps Blaming Everybody But Russia For Election Hacking - The Daily Beast #SmartNews https://t.co/KvQzjL4mHx
Newyorker2212|thedailybeast|-0.4939|0.167|0.833|0.0|RT @DerronDjjrdn: Donald Trump Keeps Blaming Everybody But Russia For Election Hacking - The Daily Beast #SmartNews https://t.co/KvQzjL4mHx
ramcatalleyetsy|_0HOUR1|-0.2235|0.079|0.921|0.0|RT @_0HOUR1: Donald Trump did not commit #Treason watch your words folks this is the President-Elect you speak of now. Especially you peopl
HelenEckard|randyprine|0.3612|0.079|0.753|0.168|"RT @randyprine: Instead of vilifying the CIA, Trump should release his taxes to prove that Russia has no incentive for helping him be elect"
Zhape|SeabreezeCheryl|-0.2808|0.172|0.71|0.118|"RT @SeabreezeCheryl: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/ufmcVURB1v via @Bipart"
Zhape|bipartisanreport|-0.2808|0.172|0.71|0.118|"RT @SeabreezeCheryl: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/ufmcVURB1v via @Bipart"
bhandarirupes18|KanakManiDixit|-0.3869|0.102|0.898|0.0|"RT @KanakManiDixit: ""Our first task in this struggle is to understand what we face.Only then can we work out what to do.""-George Monibot ht"
tlhenson823|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
LaOkieKat|asamjulian|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
LaOkieKat|twitter|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
Martina|DavidCornDC|0.8458|0.042|0.651|0.307|@DavidCornDC a very good point.But then what is trump serious about exactly We know he wants to be more wealthy and more popular? What else?
uncagedgypsy|leahmcelrath|0.0|0.0|1.0|0.0|"RT @leahmcelrath: This is a thorough compilation on @dailykos of resources regarding Putin, Dugin, Spencer, Bannon, and Trump:https://t.c"
uncagedgypsy||0.0|0.0|1.0|0.0|"RT @leahmcelrath: This is a thorough compilation on @dailykos of resources regarding Putin, Dugin, Spencer, Bannon, and Trump:https://t.c"
Mom9Ky|TheDemocrats|0.5514|0.0|0.818|0.182|RT @TheDemocrats: Are you:- A woman?- Under 26?Do you:- Have a pre-existing condition?- Live?- Breathe?Obamacare helps you. Don't le
KurtRexCooper|tomtomorrow|-0.3818|0.106|0.894|0.0|"I process Trump's cabinet picks that way.  I grieve for America at each pick, then do not think about it until the next one. @tomtomorrow"
jesse74henson|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
CHURCHLADY320|CitizensFedUp|0.2023|0.0|0.872|0.128|"RT @CitizensFedUp: Hillary could have legal right to challenge electoral college system and be next US president, says law professor https:"
tmogul_live|youtube|-0.2942|0.244|0.582|0.174|"Who Cares About Yemen's War, Trump is Person of the Year! https://t.co/xgeyIqxSRi"
MelindaThinker|SheSternly|-0.7065|0.218|0.782|0.0|"RT @SheSternly: Petition your Senators that trump is part of a proven coup by Russian forces and they know it. NO INAUGURATION, NO COOPERAT"
IntrovertRN1975|JuddLegum|0.5979|0.0|0.811|0.189|"RT @JuddLegum: 6. According to Bolton, Russians are so good at hacking they would never leave evidence that US intel could detect https://t"
IntrovertRN1975||0.5979|0.0|0.811|0.189|"RT @JuddLegum: 6. According to Bolton, Russians are so good at hacking they would never leave evidence that US intel could detect https://t"
JackieMcReath1|alexjonesshows|-0.4019|0.162|0.838|0.0|RT @alexjonesshows: Trump dismisses the CIAs claim it has evidence Russians hacked the election https://t.co/BlIQajTzOd
JackieMcReath1|alexjonespodcast|-0.4019|0.162|0.838|0.0|RT @alexjonesshows: Trump dismisses the CIAs claim it has evidence Russians hacked the election https://t.co/BlIQajTzOd
NewsBry|newsbry|0.0|0.0|1.0|0.0|"Despite scientific consensus, Trump says nobody knows if climate change isrea https://t.co/9SvBByM5wt"
lindadoherty4|kurteichenwald|0.7089|0.0|0.772|0.228|"RT @kurteichenwald: Trump says: So smart doesnt need daily intel briefings, knows more about ISIS than military, knows tax code better than"
BalanceInNature|sarahkendzior|-0.0258|0.196|0.613|0.19|RT @sarahkendzior: US Intelligence agencies fear reprisals over Russia revelations https://t.co/PP9qzrbB3s https://t.co/qwwUMIs3rV
BalanceInNature|theguardian|-0.0258|0.196|0.613|0.19|RT @sarahkendzior: US Intelligence agencies fear reprisals over Russia revelations https://t.co/PP9qzrbB3s https://t.co/qwwUMIs3rV
MarEnrile|TeenVogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
MarEnrile|teenvogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
ruthsias|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
BonnieLynn52|HAWofPA|-0.3182|0.113|0.887|0.0|@HAWofPA Trump met with Al Gore and Leo DiCaprio-he's studying this-might just be a bunch of bull for greedy politicians
bfinstock2_0|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
diamondnill1|puppymnkey|0.0|0.0|1.0|0.0|RT @puppymnkey: This one is appropriate for today. IMPEACH the TRAITOR TRUMP @speakerryan https://t.co/KXTmsGsDIx
diamondnill1|twitter|0.0|0.0|1.0|0.0|RT @puppymnkey: This one is appropriate for today. IMPEACH the TRAITOR TRUMP @speakerryan https://t.co/KXTmsGsDIx
ChicagoCro|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/X96opIoxXJ https://t.co/SpvgwkGPoS
ChicagoCro|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/X96opIoxXJ https://t.co/SpvgwkGPoS
arielvalentin|KatzOnEarth|0.4767|0.086|0.706|0.208|RT @KatzOnEarth: The Trump presidency will be dedicated to making sure everything he falsely accused Obama of doing now happens: https://t.
arielvalentin||0.4767|0.086|0.706|0.208|RT @KatzOnEarth: The Trump presidency will be dedicated to making sure everything he falsely accused Obama of doing now happens: https://t.
MariaEl26012179|EP_EEUU_24Horas|0.0|0.0|1.0|0.0|RT @EP_EEUU_24Horas: Billete parejo! El gabinete de Trump colmado de millonarios https://t.co/XXiaCiA4kN https://t.co/kbNdPuE168
MariaEl26012179|epmundo|0.0|0.0|1.0|0.0|RT @EP_EEUU_24Horas: Billete parejo! El gabinete de Trump colmado de millonarios https://t.co/XXiaCiA4kN https://t.co/kbNdPuE168
GoodHumorGrl|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
zmain1|Joyce_Karam|-0.8176|0.309|0.691|0.0|RT @Joyce_Karam: There's an attack on Church in Egypt;Terror in Istanbul; ISIS took Palmyra; CIA alarm on Russia.But #Trump is attacking NB
sud_vijay|kurteichenwald|0.7089|0.0|0.772|0.228|"RT @kurteichenwald: Trump says: So smart doesnt need daily intel briefings, knows more about ISIS than military, knows tax code better than"
Daniel7964|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
remmkm|Adenovir|-0.8658|0.386|0.614|0.0|"RT @Adenovir: Carl Bernstein, who broke the Watergate scandal that led to Nixon's resignation, said that Nixon's lies were nothing compared"
nancy73gg|LindaSuhler|0.0|0.0|1.0|0.0|"RT @LindaSuhler: #PEOTUS Donald J. Trump #ThankYouTour2016 #FloridaOrlando, FLFRIDAY 7 PM ET#MAGA #AmericaFirstRegis:https://t.co"
nancy73gg|t|0.0|0.0|1.0|0.0|"RT @LindaSuhler: #PEOTUS Donald J. Trump #ThankYouTour2016 #FloridaOrlando, FLFRIDAY 7 PM ET#MAGA #AmericaFirstRegis:https://t.co"
meaghanwebster|nytimes|0.0|0.0|1.0|0.0|"RT @nytimes: Rex Tillerson, the Exxon Mobil chief with ties to Putin, is expected to be Trump's pick for secretary of state https://t.co/7A"
meaghanwebster|t|0.0|0.0|1.0|0.0|"RT @nytimes: Rex Tillerson, the Exxon Mobil chief with ties to Putin, is expected to be Trump's pick for secretary of state https://t.co/7A"
ReclaimDawgs|TeaPartyCore|0.743|0.0|0.687|0.313|RT @TeaPartyCore: values and principles of #TeaParty movement r finally gaining the top seat of power in the White Househttps://t.co/QMDfn
drv4posgrowth|JimmyBear2|-0.1779|0.188|0.663|0.149|"RT @JimmyBear2: POLITIFACT: Trump Is Lying, Russia DID Swing Election In His Favor - https://t.co/10wfG8wcui"
drv4posgrowth|occupydemocrats|-0.1779|0.188|0.663|0.149|"RT @JimmyBear2: POLITIFACT: Trump Is Lying, Russia DID Swing Election In His Favor - https://t.co/10wfG8wcui"
PedroCo16889625|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
kehindekolawole|KatyTurNBC|0.4215|0.0|0.823|0.177|@KatyTurNBC when are u writing a book sharing your experience on the campaign trail with Trump ?
hypnocoach183|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
sa_solomon|washingtonpost|-0.1531|0.106|0.817|0.077|"After asking Who believes in global warming? &amp; soliciting a show of hands, Trump concluded no one did. #IdiotinChief https://t.co/00NrHzj787"
Maxzen2004|TheTrumpLady|0.4184|0.133|0.625|0.242|"RT @TheTrumpLady: Wow! Unbelievable! #Ryan Working With Trump on Wall, Deport Criminal Illegals, Extreme Vetting, School Choice, etc. https"
4EverJohnnyBoy|NancyLeeGrahn|-0.1779|0.218|0.627|0.155|@NancyLeeGrahn SO rad see you in my notifications. Love Alexis &amp; need #GeneralHospital to distract from insanity of #Trump #TrumpTransition.
SFH26|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
B_H_Fan4Evr|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
an_janes|divinity254|0.4588|0.0|0.864|0.136|RT @divinity254: GM @AlohaMsLonesome Trump only cares about himself &amp; lining his pockets. Troops? He doesn't even attend daily briefings @
uramkmf4|dailykos|0.0|0.0|1.0|0.0|Rachel Maddow: Poll reveals Trump voters live in alternate state of reality https://t.co/quD1b4tfr5
1549321s|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: US Senators letter to Senate leaders-investigate Trump for Russian espionage#cnn #msnbc #AMJoy #cnnsotu #thiswee
BelkissObadia|TeaPainUSA|-0.0516|0.101|0.804|0.094|RT @TeaPainUSA: Now we see clearly why Trump wants to abandon NATO &amp; give Putin the green light to rebuild the old Soviet empire. #RedDon #
llarks|ckilpatrick|0.2042|0.12|0.693|0.186|RT @ckilpatrick: Trump will not be defeated by outrage. He'll be defeated by (socialist) Left populist politics. We should be most concerne
GoodwinHH6|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
MarieFrRenaud|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
dal4kids|SPNlocal|0.0|0.0|1.0|0.0|@SPNlocal @RealBenCarson @ALLNCom @realDonaldTrump @Trump @mikepence @ArcLight_Cares @choice_renovate  https://t.co/ODy53pI0Qo
dal4kids|linkedin|0.0|0.0|1.0|0.0|@SPNlocal @RealBenCarson @ALLNCom @realDonaldTrump @Trump @mikepence @ArcLight_Cares @choice_renovate  https://t.co/ODy53pI0Qo
ar1511c|JSavoly|-0.0258|0.114|0.778|0.108|RT @JSavoly: Top Republicans Just Demanded An Investigation Into Russia's Pro-Trump Interference #StollenElection #ComradeTrump  https://t.
ar1511c||-0.0258|0.114|0.778|0.108|RT @JSavoly: Top Republicans Just Demanded An Investigation Into Russia's Pro-Trump Interference #StollenElection #ComradeTrump  https://t.
roznewz|thehill|0.0|0.0|1.0|0.0|RT @thehill: Trump goes after NBC news in tweethttps://t.co/32I8myfDsw https://t.co/vj13vixfUJ
roznewz|twitter|0.0|0.0|1.0|0.0|RT @thehill: Trump goes after NBC news in tweethttps://t.co/32I8myfDsw https://t.co/vj13vixfUJ
JackEddieFoster|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
ThomasJankow|squad19mpls|0.6705|0.0|0.703|0.297|"RT @squad19mpls: I'm pretty sure Trump is the first self-serving asshole to be president, ever."
MLorance|RepAdamSchiff|-0.34|0.118|0.882|0.0|RT @RepAdamSchiff: There's overwhelming evidence of Russian hacking of our elections. By denying it Trump has essentially become a propagan
sosarcatstic|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
sosarcatstic|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
mikehaddad|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
mikehaddad|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
Apipwhisperer|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
Apipwhisperer||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
paulrlanni|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
paulrlanni|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
TheJakeMassaro|DRUDGE_REPORT|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: 'FACTS ARE THERE' https://t.co/lIkm59zJrx
TheJakeMassaro|cbsnews|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: 'FACTS ARE THERE' https://t.co/lIkm59zJrx
SuzanneinLGB|Khanoisseur|-0.4588|0.15|0.85|0.0|RT @Khanoisseur: 2 reasons for trump rejecting daily intel briefings:1. Plausible deniability2. Busy making side deal$$ for himself @mrp
nia4_trump|mikandynothem|0.7845|0.0|0.717|0.283|RT @mikandynothem: John Kenedy wins last seat in landslide for Senate giving #GOP 52-48 majority. The cherry on the top of a Republican Rev
PaytonBennett5|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
PaytonBennett5|thegatewaypundit|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
AlexTheGreatzz|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
saraewelch1|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
saraewelch1||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
pabl_ohhh|AdamSmith_usa|0.0|0.0|1.0|0.0|RT @AdamSmith_usa: This fleece has more experience than Donald Trump. https://t.co/USGojcf5lX
pabl_ohhh|twitter|0.0|0.0|1.0|0.0|RT @AdamSmith_usa: This fleece has more experience than Donald Trump. https://t.co/USGojcf5lX
Paidsubscriber|burnaby1953|0.4939|0.127|0.615|0.258|RT @burnaby1953: Dan Rather Just Called Out Fake Patriots Who Support Trumps Putin Romance In Viral Post - https://t.co/2tJcaY0PP8
Paidsubscriber|occupydemocrats|0.4939|0.127|0.615|0.258|RT @burnaby1953: Dan Rather Just Called Out Fake Patriots Who Support Trumps Putin Romance In Viral Post - https://t.co/2tJcaY0PP8
rdnktk|tonyschwartz|-0.296|0.091|0.909|0.0|RT @tonyschwartz: I don't believe anything Donald Trump says. Not one word. It is all manipulation and mind games all the time. (Same for K
NadiaGladysM|Toure|0.6647|0.113|0.532|0.355|RT @Toure: Trump says he doesnt need intelligence briefings because Im a smart person. God save us.
Tech_Stuff_Go|washingtonpost|0.0|0.0|1.0|0.0|Six Of Trump's Cabinet Appointees Gave Almost $12 Million To Trump's Campaign https://t.co/JfASExo8IS
hawaiianlove68|tribelaw|-0.5106|0.125|0.875|0.0|RT @tribelaw: But mounting public outrage at Trump's benefiting his family business at the expense of U.S. working men and women will do hi
DerpyPhlllip|DrJenGunter|-0.5994|0.205|0.795|0.0|RT @DrJenGunter: If Trump is right and there was no Russian interference what does he have to lose from an investigation?
KimbaGross|Mama3Cubs|0.5719|0.0|0.778|0.222|"RT @Mama3Cubs: @Astorix23 @Bow2kaos The only thing ""foreign"" to Donald Trump is success: https://t.co/X53DPHtPZu"
KimbaGross|twitter|0.5719|0.0|0.778|0.222|"RT @Mama3Cubs: @Astorix23 @Bow2kaos The only thing ""foreign"" to Donald Trump is success: https://t.co/X53DPHtPZu"
sweetteatime55|WilliamCohan|-0.25|0.124|0.796|0.08|Trump cheats while playing golf @WilliamCohan Author of Money and Power House of Cards The Last Tycoon speaks on https://t.co/2BmYJVEDVG
sweetteatime55|twitter|-0.25|0.124|0.796|0.08|Trump cheats while playing golf @WilliamCohan Author of Money and Power House of Cards The Last Tycoon speaks on https://t.co/2BmYJVEDVG
SonofCarnelian|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
blueinthesouth|MarkHarrisNYC|-0.8555|0.331|0.669|0.0|RT @MarkHarrisNYC: Those briefings scare Trump--they're full of info he doesn't know and can't hold onto. And being scared angers him.  htt
chicagogrrrl|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
chicagogrrrl|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
RemiPerry|CaptainsLog2016|0.0|0.119|0.72|0.161|RT @CaptainsLog2016: Donald Trump said this word for wordOn national television&amp; now denies believing in any chance of Russia playing a
NorthernPikeFly|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
ElaineLafon|NBCNews|0.0516|0.145|0.661|0.194|RT @NBCNews: A slap in the face. That's how intelligence agencies see Trump's rejection of findings on Russia https://t.co/k6QZxwjtem https
ElaineLafon|nbcnews|0.0516|0.145|0.661|0.194|RT @NBCNews: A slap in the face. That's how intelligence agencies see Trump's rejection of findings on Russia https://t.co/k6QZxwjtem https
jyester55|KeithOlbermann|0.3818|0.0|0.902|0.098|"RT @KeithOlbermann: HOW could Russians run coup to elect the disloyal Trump? From 12/2: when they try to hack YOU, the answer is clear: htt"
KPHennosy|tribelaw|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
KPHennosy|twitter|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
Superjew75|twitter|0.5106|0.097|0.686|0.217|This thread is a fantastic analysis of how we got to Russia giving us President Trump &amp; him ignoring CIA/FBI &amp; obvi https://t.co/W3RUBoIxbE
kikidasu1|BruceBartlett|0.5106|0.0|0.82|0.18|RT @BruceBartlett: Strong evidence that FBI Director Comey delivered the White House to Trump. https://t.co/k5q4Sn56bt https://t.co/WCr5kvF
kikidasu1|election|0.5106|0.0|0.82|0.18|RT @BruceBartlett: Strong evidence that FBI Director Comey delivered the White House to Trump. https://t.co/k5q4Sn56bt https://t.co/WCr5kvF
philippberner|recode|0.0|0.0|1.0|0.0|"What Trump said about Apple, Alphabet and Facebook  the tech companies hes meeting next week - Recode https://t.co/7M4T0aliNU"
tammy_wesa|Khanoisseur|0.0772|0.0|0.925|0.075|RT @Khanoisseur: He actually gave this as an excuse for skipping daily ntelligence briefings https://t.co/xG4TtdK7QB @Green_Footballs @kurt
tammy_wesa|washingtonpost|0.0772|0.0|0.925|0.075|RT @Khanoisseur: He actually gave this as an excuse for skipping daily ntelligence briefings https://t.co/xG4TtdK7QB @Green_Footballs @kurt
LKuehn4|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
KatEdmiston|gollum1419_g|0.0|0.0|1.0|0.0|RT @gollum1419_g: Possible Trump Appointee Scrubs Facebook Post Fantasizing About Exterminating Muslims https://t.co/m3W7xL65AK #Resist #Tr
KatEdmiston|rawstory|0.0|0.0|1.0|0.0|RT @gollum1419_g: Possible Trump Appointee Scrubs Facebook Post Fantasizing About Exterminating Muslims https://t.co/m3W7xL65AK #Resist #Tr
fhs_PACE|yearbook_falcon|0.4404|0.0|0.838|0.162|"@yearbook_falcon &amp; @aggresivespice are interviewing trump/bernie/clinton supporters, &amp; our gen meet is wed, so come thru "
GagaDelRey25|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
sciencemilkcow|Joyce_Karam|0.0|0.0|1.0|0.0|"RT @Joyce_Karam: Not one tweet or word on Egypt or Turkey from Trump. If those intel briefings are repetitive/boring, how about start with"
johnobmickel|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
IntrovertRN1975|JuddLegum|-0.3612|0.111|0.889|0.0|"RT @JuddLegum: 5. Bolton's evidence of this is that the CIA found evidence of Russian involvement, which he finds suspicious https://t.co/o"
IntrovertRN1975|twitter|-0.3612|0.111|0.889|0.0|"RT @JuddLegum: 5. Bolton's evidence of this is that the CIA found evidence of Russian involvement, which he finds suspicious https://t.co/o"
PriyankaVakil|BrookingsInst|0.0|0.0|1.0|0.0|RT @BrookingsInst: 46% of Americans think Obama should take action on Israel-Palestine before leaving office https://t.co/pr01irnpBj https:
PriyankaVakil|brookings|0.0|0.0|1.0|0.0|RT @BrookingsInst: 46% of Americans think Obama should take action on Israel-Palestine before leaving office https://t.co/pr01irnpBj https:
CNNedition|cnn|0.0|0.0|1.0|0.0|Trump: 'Nobody really knows' if climate change is real https://t.co/Z6Py9VoS1W
TurnTNBlue|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
trumpfnd|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
Wyohawk|DailyCaller|-0.7603|0.361|0.459|0.18|"RT @DailyCaller: Kellyanne Conway, After Getting Death Threats, EPICALLY DESTROYS People Who Just Cant Admit Trump Won [VIDEO] https://t"
Wyohawk||-0.7603|0.361|0.459|0.18|"RT @DailyCaller: Kellyanne Conway, After Getting Death Threats, EPICALLY DESTROYS People Who Just Cant Admit Trump Won [VIDEO] https://t"
IqbalSharifBiru|twitter|0.3818|0.0|0.874|0.126|"Dear Fox News,Donald J.Trump is the elected President of U.S.And it should duly be respected.Please see my Facebook https://t.co/Niq4zpxqPR"
querderai|fperez_org|-0.128|0.174|0.711|0.115|"RT @fperez_org: The US did stop the McCarthy era, will it stop its modern renaissance? Good perspective from Adorno et al.:https://t.co/0F"
querderai|t|-0.128|0.174|0.711|0.115|"RT @fperez_org: The US did stop the McCarthy era, will it stop its modern renaissance? Good perspective from Adorno et al.:https://t.co/0F"
DavidPoland|SeanMcElwee|0.6249|0.0|0.796|0.204|"RT @SeanMcElwee: Trump gave cabinet positions to 6 major donors, which is unprecedented. Great reporting from @mateagold. https://t.co/2w4v"
DavidPoland|t|0.6249|0.0|0.796|0.204|"RT @SeanMcElwee: Trump gave cabinet positions to 6 major donors, which is unprecedented. Great reporting from @mateagold. https://t.co/2w4v"
ltowsonhester|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
Presley48R|TeamTrumpCO|0.6027|0.0|0.781|0.219|RT @TeamTrumpCO: now 5K followers THANKS! Began in spring16.Tweeted 4 #Leave &amp; #Brexit &amp; #MAGA3X&amp; #Trump.#antieu#antiglobalism#AmericaFi
madmatt015|realDonaldTrump|-0.5619|0.25|0.647|0.103|"@realDonaldTrump @NBCNightlyNews @CNN Just read Trump' tweets- So biased, inaccurate &amp; bad, point after point. Can't get much worse!"
John72115John|politico|-0.8713|0.397|0.603|0.0|"@politico @SpeakerRyan IF RYAN HAD A SCROTUM, MAYBE HE'D STEP UP N EXPOSE TRUMP! NAH! TOO MUCH BITCH IN HIM!"
TootiePalmer|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
JHSaunders|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Trump eyes TAIWAN for luxury home projects-he does biz there#cnn #msnbc #amjoy #maddow #fridayfeeling https://t.
JHSaunders||0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Trump eyes TAIWAN for luxury home projects-he does biz there#cnn #msnbc #amjoy #maddow #fridayfeeling https://t.
PaulJAndrew|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
heresursign_1|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
babysgramma|rtoberl|0.2732|0.0|0.87|0.13|RT @rtoberl: Supposedly tolerant NYC is making the Trump kids' lives 'horrible' https://t.co/hbxgESyvc6 via @nypost
babysgramma|linkis|0.2732|0.0|0.87|0.13|RT @rtoberl: Supposedly tolerant NYC is making the Trump kids' lives 'horrible' https://t.co/hbxgESyvc6 via @nypost
zackola|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
zackola|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
FlavioCastroSay|Forbes|0.0|0.0|1.0|0.0|RT @Forbes: Take a look inside Trump's $100 million private jet: https://t.co/CfrvKeExGp https://t.co/Ar3DfhnLOH
FlavioCastroSay|forbes|0.0|0.0|1.0|0.0|RT @Forbes: Take a look inside Trump's $100 million private jet: https://t.co/CfrvKeExGp https://t.co/Ar3DfhnLOH
burmoll|Anncostanza1|0.902|0.0|0.598|0.402|RT @Anncostanza1: Trump Knocked it out of the Park with Secretary of Defense General MadDogMattis Awesome! Respect our Troops Respect US Fl
NatashaDargan|JoshButler|0.0|0.0|1.0|0.0|"RT @JoshButler: The New York Times piece on Australia's refugee policy is blistering. Dutton is our ""little Trump""  https://t.co/hvwnJ7XV7O"
NatashaDargan|mobile|0.0|0.0|1.0|0.0|"RT @JoshButler: The New York Times piece on Australia's refugee policy is blistering. Dutton is our ""little Trump""  https://t.co/hvwnJ7XV7O"
JackieMcReath1|LVNancy|0.5719|0.0|0.791|0.209|"RT @LVNancy: #RussianHackers IF sore-Loser, Hillary had won, would we be having this conversation?#SundayMorning #TRUMP#AmericaFirst"
anobscureartist|EdSkipper|0.765|0.0|0.752|0.248|RT @EdSkipper: Wisely most of Europe wanted a Clinton win. But they didn't meddle. #RussianHacking did. Comey knew. US Intel knows. Did Tru
nancy73gg|LindaSuhler|0.0|0.0|1.0|0.0|"RT @LindaSuhler: #PEOTUS Donald J. Trump #ThankYouTour2016 #AlabamaMobile, ALSaturday, 3 PM CT#MAGA #AmericaFirstRegis:https://t."
nancy73gg||0.0|0.0|1.0|0.0|"RT @LindaSuhler: #PEOTUS Donald J. Trump #ThankYouTour2016 #AlabamaMobile, ALSaturday, 3 PM CT#MAGA #AmericaFirstRegis:https://t."
NoMoreElites|jimlibertarian|0.0|0.0|1.0|0.0|"RT @jimlibertarian: Jan 20th of 2017 will mark the beginning of a new era,Donald Trump will B our 45th POTUS https://t.co/3WMUu48sUn htt"
NoMoreElites|i|0.0|0.0|1.0|0.0|"RT @jimlibertarian: Jan 20th of 2017 will mark the beginning of a new era,Donald Trump will B our 45th POTUS https://t.co/3WMUu48sUn htt"
masonbo|gatewaypundit|0.128|0.111|0.754|0.136|RT @gatewaypundit: FBI Investigation Refutes CIA=&gt; Theres No Evidence Russia Tried to Help Trump https://t.co/7epYPdIaUF via @gatewaypundit
masonbo|thegatewaypundit|0.128|0.111|0.754|0.136|RT @gatewaypundit: FBI Investigation Refutes CIA=&gt; Theres No Evidence Russia Tried to Help Trump https://t.co/7epYPdIaUF via @gatewaypundit
noahastevens|twitter|0.0|0.0|1.0|0.0|this should get the Trump folks riled up: https://t.co/MTvTTyWOtV
VagabondWahine|twitter|-0.6249|0.231|0.769|0.0|"Either Trump knew Russia was manipulating elections, which makes him  corrupt, or he let himself be manipulated, wh https://t.co/tWRR0dn82c"
KRCSmith62|ThePCJF|0.4404|0.062|0.793|0.145|"RT @ThePCJF: National Park Service ""has done a massive land grab"" inhibiting free speech rights on Inauguration Day via @Reuters https://t."
KRCSmith62||0.4404|0.062|0.793|0.145|"RT @ThePCJF: National Park Service ""has done a massive land grab"" inhibiting free speech rights on Inauguration Day via @Reuters https://t."
HMKohnlein|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
SheSternly|twitter|-0.7829|0.293|0.707|0.0|trump has no more validity w/his fantasy of running our country for Russia. Do not help him normalize this. STOP TH https://t.co/zOEuXR458t
roqchrisy|LouDobbs|0.0|0.0|1.0|0.0|RT @LouDobbs: The New Boss is the New Boss!  #MAGA #AmericaFirst #Trump #Dobbs https://t.co/zrHGqeKI7B
roqchrisy|twitter|0.0|0.0|1.0|0.0|RT @LouDobbs: The New Boss is the New Boss!  #MAGA #AmericaFirst #Trump #Dobbs https://t.co/zrHGqeKI7B
trumpfnd|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
angxlthenerd|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
522tim|Poynter|-0.5267|0.195|0.805|0.0|"RT @Poynter: Donald Trump's real threat to the press? The Espionage Act, not libel laws.https://t.co/3vVmgWQ1Je"
Seacretsoc1|ExportedFromMI|-0.0772|0.142|0.728|0.13|RT @ExportedFromMI: @JuddLegum Where is Chief Justice John Roberts? Borderline treasonous activity from the Trump team &amp; only a few GOP con
RichandGod|twitter|-0.0772|0.154|0.71|0.136|Donald Trump told us the truth that's why he's president Hillary lied consistently https://t.co/hQAp5JKWMC
ramzpaul|Communism_Kills|0.5719|0.0|0.829|0.171|"RT @Communism_Kills: Here is a perfect example of #fakenews: a story about a tweet and my ""sexist"" reply to the tweet. https://t.co/yh5MHQj"
ramzpaul|t|0.5719|0.0|0.829|0.171|"RT @Communism_Kills: Here is a perfect example of #fakenews: a story about a tweet and my ""sexist"" reply to the tweet. https://t.co/yh5MHQj"
croneclone|davidsirota|0.0|0.0|1.0|0.0|RT @davidsirota: REVEALED: Docs show Exxon lobbied the State Dept on Russia &amp; Iran sanctions - now Exxon's CEO may run the State Dept https
LaVerneWright13|starfirst|0.4404|0.0|0.854|0.146|RT @starfirst: Fox contributor Judy Miller calls investigation of Russian hacking Obamas tar baby gift to Trump https://t.co/CpWQr2Eepb
LaVerneWright13|rawstory|0.4404|0.0|0.854|0.146|RT @starfirst: Fox contributor Judy Miller calls investigation of Russian hacking Obamas tar baby gift to Trump https://t.co/CpWQr2Eepb
Willie_Jacobsz|greenhousenyt|0.0|0.0|1.0|0.0|RT @greenhousenyt: NYT EditorialTrump should lead call for a thorough investigation. It's only way to remove cloud from his presidency htt
ScorpiusDragon|rstevens|0.3818|0.105|0.673|0.222|"RT @rstevens: Hate to admit it, but I support Trumps choice of Cigarette Smoking Man for Surgeon General https://t.co/QDvLTsca85"
ScorpiusDragon|twitter|0.3818|0.105|0.673|0.222|"RT @rstevens: Hate to admit it, but I support Trumps choice of Cigarette Smoking Man for Surgeon General https://t.co/QDvLTsca85"
sampson_elaine|carlreiner|-0.34|0.208|0.66|0.132|"RT @carlreiner: As elated as I was about seeing Dick Van Dyke Show In color tonite, that's how depressed I am about Trump's choices for U.S"
FrankJannuzi|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/jWaCzABizw https://t.co/mD7GzZCYaf
FrankJannuzi|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/jWaCzABizw https://t.co/mD7GzZCYaf
randyshort|realalexjones|-0.5719|0.222|0.778|0.0|STUDY: 77 percent of Trumps general election news coverage was negative https://t.co/JjLrTGrGrB via @realalexjones
randyshort|infowars|-0.5719|0.222|0.778|0.0|STUDY: 77 percent of Trumps general election news coverage was negative https://t.co/JjLrTGrGrB via @realalexjones
redhead4645|cala_1111|0.2677|0.136|0.639|0.225|"RT @cala_1111: OPINION : Its not Trump thats a ""Danger to America,"" It's Talking Heads Like Hateful Megyn Kelly https://t.co/E0vasSxlNN"
redhead4645|truthfeed|0.2677|0.136|0.639|0.225|"RT @cala_1111: OPINION : Its not Trump thats a ""Danger to America,"" It's Talking Heads Like Hateful Megyn Kelly https://t.co/E0vasSxlNN"
stanthemanchan|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
AkSporting76|Khanoisseur|0.5859|0.0|0.84|0.16|"RT @Khanoisseur: One of the most underreported stories: How Russian money powered Trump's financial comeback, helped him win the White Hous"
reachout2015B|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
HansAlbright|BernieSanders|-0.1531|0.122|0.778|0.1|RT @BernieSanders: Donald Trump is a pathological liar.  We need the help of the American people to build a movement of millions who are fo
laughinghyena13|jayrosen_nyu|-0.2144|0.074|0.926|0.0|"RT @jayrosen_nyu: 19/ The problem is not at the level ""how to cover Trump,"" but how to recover conditions in which anything journalists do"
MikeHighley1|Mike_Beacham|0.0|0.0|1.0|0.0|RT @Mike_Beacham: Kellyanne Conway: Tillerson is part of the 'Trump effect' https://t.co/m81apFUVyd
MikeHighley1|video|0.0|0.0|1.0|0.0|RT @Mike_Beacham: Kellyanne Conway: Tillerson is part of the 'Trump effect' https://t.co/m81apFUVyd
HASSIA|RadioFreeTom|0.4767|0.0|0.876|0.124|"RT @RadioFreeTom: If HRC chose a SecState who ran an oil giant and got a medal from Putin, the GOPers defending Trump would re-convene the"
MomoAdalois|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
IntrovertRN1975|JuddLegum|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
IntrovertRN1975|t|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
FimusTauri|bbc5live|0.0|0.0|1.0|0.0|"@bbc5live Just to be topical, does Neville cringe as much as I at Trump's use of ""bigly""?"
Dbiggs1007Donna|TomthunkitsMind|-0.743|0.249|0.671|0.08|RT @TomthunkitsMind: You Can Tell By Trump's Staff Picks That We Are Going To War Within 2 Years. It's A War Cabinet. Get Ready For A Possi
djsandwiches|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
MrShellBlog|CyberHitchhiker|0.0|0.0|1.0|0.0|RT @CyberHitchhiker: Donald Trump on Russian hacking: 'I don't believe it' - https://t.co/pFVmqxU4oB https://t.co/jg2JpQzoW5 #Hacking #News
MrShellBlog|myfox8|0.0|0.0|1.0|0.0|RT @CyberHitchhiker: Donald Trump on Russian hacking: 'I don't believe it' - https://t.co/pFVmqxU4oB https://t.co/jg2JpQzoW5 #Hacking #News
lizfitz123|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
lizfitz123|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
bobgerbasi|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
bobgerbasi|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
Reggiebub|mikeallen|0.2006|0.095|0.776|0.129|"RT @mikeallen: .@jimrutenberg column salutes @jaketapper: ""If only such moments could stop being so special and start being normal"" https:/"
Reggiebub||0.2006|0.095|0.776|0.129|"RT @mikeallen: .@jimrutenberg column salutes @jaketapper: ""If only such moments could stop being so special and start being normal"" https:/"
Politolizer|politics|0.4019|0.0|0.828|0.172|Wash Post: Trumps Election Stole My Desire to Look for a Partner - Breitbart... https://t.co/uKdp869VA3 https://t.co/g5DL6RpXP3
SDPacificBeach|OANN|-0.6249|0.159|0.841|0.0|"@OANN Of course the Russkies hacked both DNC &amp; RNC &amp; of course, they wanted DT, &amp; of course they now have a lot of dirt on RNC too. Ha#Trump"
Michell66010778|joshrogin|0.1027|0.098|0.784|0.118|RT @joshrogin: .@RepAdamSchiff points out that Trump is basically giving Russia endless propaganda material at this point. @MeetThePress
addykateglen|agearan|0.631|0.0|0.813|0.187|RT @agearan: The statement does not mention Trump but still. Intelligence professionals aren't given to making such statements. https://t.c
addykateglen||0.631|0.0|0.813|0.187|RT @agearan: The statement does not mention Trump but still. Intelligence professionals aren't given to making such statements. https://t.c
khuja2006|Reuters|0.0|0.0|1.0|0.0|RT @Reuters: McCain to Trump on Russian hacking: 'The facts are there' - CBS https://t.co/QoesspVeoq https://t.co/pP6xj54U5Q
khuja2006|reuters|0.0|0.0|1.0|0.0|RT @Reuters: McCain to Trump on Russian hacking: 'The facts are there' - CBS https://t.co/QoesspVeoq https://t.co/pP6xj54U5Q
SharonS72105601|LouDobbs|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
SharonS72105601|theconservativetreehouse|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
dogfriendlydude|SenSanders|0.4767|0.08|0.691|0.229|"RT @SenSanders: I challenge Mr. Trump to tell the American people he'll keep his promises and veto cuts to Social Security, Medicare and Me"
soozanderson4|MikeBates|0.4019|0.0|0.803|0.197|"RT @MikeBates: Unnecessary for such a smart person. He watches ""the shows.""  https://t.co/QrSvis4mYr"
soozanderson4|businessinsider|0.4019|0.0|0.803|0.197|"RT @MikeBates: Unnecessary for such a smart person. He watches ""the shows.""  https://t.co/QrSvis4mYr"
stilllwithher|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
stilllwithher|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
Deplorable80210|laurenduca|-0.3535|0.127|0.873|0.0|@laurenduca @TeenVogue's journalism is just more #FAKENEWS ... Missed a VERY BIG PROOF GAP on the Russia hacking https://t.co/WfhzF8fo03
Deplorable80210|cnn|-0.3535|0.127|0.873|0.0|@laurenduca @TeenVogue's journalism is just more #FAKENEWS ... Missed a VERY BIG PROOF GAP on the Russia hacking https://t.co/WfhzF8fo03
djpriller|dayvarelat|0.128|0.0|0.914|0.086|RT @dayvarelat: Exclusive  First Day of Trumps Presidency: President-Elect Highlights Sacrifice of Americas Armed Forces at https://t
djpriller||0.128|0.0|0.914|0.086|RT @dayvarelat: Exclusive  First Day of Trumps Presidency: President-Elect Highlights Sacrifice of Americas Armed Forces at https://t
lsuagain|PSheritaakkloh|-0.6199|0.238|0.762|0.0|"@PSheritaakkloh @JhoniiAlmeida If you hate Trump, why are you following his tweets? Troll much?"
sublett_pamelia|kurteichenwald|-0.5423|0.176|0.824|0.0|"RT @kurteichenwald: Fox/Cheney went nuts when found out Obama got intel briefings in writing, rather than read to him. But Trump no briefin"
Apipwhisperer|FoxNews|-0.1779|0.124|0.876|0.0|RT @FoxNews: .@JudgeJeanine Slams Obama: 'Why Are You Obsessed With Russia?' https://t.co/96TVMVqFc9 https://t.co/WkwW8sYfbg
Apipwhisperer|insider|-0.1779|0.124|0.876|0.0|RT @FoxNews: .@JudgeJeanine Slams Obama: 'Why Are You Obsessed With Russia?' https://t.co/96TVMVqFc9 https://t.co/WkwW8sYfbg
AskMrPickles|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
cosmicsource|CollectiveEvol|0.0|0.0|1.0|0.0|"@CollectiveEvol the Trump clip from the Simpsons isn't from 2000, it came out after the real footage https://t.co/eareWKgzzd"
cosmicsource|youtube|0.0|0.0|1.0|0.0|"@CollectiveEvol the Trump clip from the Simpsons isn't from 2000, it came out after the real footage https://t.co/eareWKgzzd"
Traveljunkie213|frankrichny|-0.1603|0.064|0.936|0.0|"RT @frankrichny: By holding back RNC emails, Putin didn't just help install Trump in White House but has means to blackmail GOP to do his b"
TurnTNBlue|TheDemocrats|0.5514|0.0|0.818|0.182|RT @TheDemocrats: Are you:- A woman?- Under 26?Do you:- Have a pre-existing condition?- Live?- Breathe?Obamacare helps you. Don't le
DocDonDJ|AntTheIcon|0.4515|0.141|0.617|0.242|RT @AntTheIcon: worst 2 teams? 49ers with a BLM QB and the BROWNS. best record? the AMERICAN conference PATRIOTS whose QB publicly supports
LindaWestbroo11|seankent|0.9179|0.0|0.536|0.464|"RT @seankent: Trump voters, does this seem like a legit reason for skipping intelligence briefings? Does it inspire confidence?   https://t"
LindaWestbroo11||0.9179|0.0|0.536|0.464|"RT @seankent: Trump voters, does this seem like a legit reason for skipping intelligence briefings? Does it inspire confidence?   https://t"
hypnocoach183|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
MarianMme16513|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
MarianMme16513|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
cyber_gr1zzly|buzz|-0.7269|0.307|0.693|0.0|RT @buzz: When even the foreign power manipulating you is shocked at your party's lack of principle. https://t.co/4erdcrGxSk https://t.co/8
cyber_gr1zzly|newsweek|-0.7269|0.307|0.693|0.0|RT @buzz: When even the foreign power manipulating you is shocked at your party's lack of principle. https://t.co/4erdcrGxSk https://t.co/8
going2left|NancyErvin4|0.2057|0.0|0.927|0.073|"RT @NancyErvin4: GOP in collusion with trump &amp; Russia. Knew of trump allegiance to Russia, not USA. Blocked all attempts to get to truth=ta"
surfgranma|SwissTriple_M|0.0|0.0|1.0|0.0|RT @SwissTriple_M: That is #insidertrading if he told Baer Sterns 2 buy stock based on inside information on Bally. #marthastewart did her
KeenaGreene|HuffPostPol|-0.8354|0.343|0.657|0.0|"SMH ths mf is dumb af Trump says he doesn't need a daily intelligence briefing because he's ""smart"" https://t.co/Mixp0OGpwL via @HuffPostPol"
KeenaGreene|huffingtonpost|-0.8354|0.343|0.657|0.0|"SMH ths mf is dumb af Trump says he doesn't need a daily intelligence briefing because he's ""smart"" https://t.co/Mixp0OGpwL via @HuffPostPol"
daxis_gaming|RamonaCallender|-0.1027|0.08|0.92|0.0|@RamonaCallender oh also many will try to get trump to pay for it all as he should
soytome|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soytome|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
GayRainey1|itsbrycegreene|0.1759|0.147|0.678|0.175|@itsbrycegreene @RogerJStoneJr @realDonaldTrump @YouTube I don't see how anyone could hate Mr. Trump. He is doing great things for America!
JCupcakeee|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
soycalama|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soycalama|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyvaldiviacl|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyvaldiviacl|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyvalparaiso|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyvalparaiso|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
Bilmartighan|Nate_Cohn|0.1531|0.121|0.738|0.141|RT @Nate_Cohn: I guess the Trump-Bolton case is that there were 2m illegal votes and a CIA false flag op in one of the greatest victories i
soyarica|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyarica|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soycopiapo|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soycopiapo|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soytalcahuano|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soytalcahuano|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyquillota|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyquillota|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyiquique|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyiquique|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soysanantonio|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soysanantonio|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soypuertomontt|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soypuertomontt|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyconcepcion|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyconcepcion|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyosorno|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyosorno|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soychillan|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soychillan|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soychiloe|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soychiloe|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyarauco|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyarauco|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyantofagasta|soychilecl|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
soyantofagasta|soychile|0.0|0.0|1.0|0.0|"RT @soychilecl: Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
NonaHarman|HamiltonElector|-0.296|0.099|0.901|0.0|RT @HamiltonElector: We've crossed the threshold. There is no going back. Trump must never become POTUS. RT to let #hamiltonelectors know y
corgiman3|JohnWDean|-0.6597|0.188|0.76|0.052|"RT @JohnWDean: Notwithstanding Trump's efforts to kill this, there are a few real Americans in the US Senate who want answers: https://t.co"
corgiman3|t|-0.6597|0.188|0.76|0.052|"RT @JohnWDean: Notwithstanding Trump's efforts to kill this, there are a few real Americans in the US Senate who want answers: https://t.co"
AnitaBalch|actionnetwork|0.3595|0.0|0.865|0.135|I'm mobilizing to #StopTrump and #DefendDemocracy at my state capitol on #dec19. Join us! RSVP here: https://t.co/lGLAARd025
BrianAnthonyMc|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
rob_fulwell|nebraskamlc|0.0|0.0|1.0|0.0|@nebraskamlc Well... https://t.co/V9lCwX6heY
rob_fulwell|cnn|0.0|0.0|1.0|0.0|@nebraskamlc Well... https://t.co/V9lCwX6heY
WhosFibbing|LouDobbs|-0.6597|0.221|0.779|0.0|RT @LouDobbs: The Ignorance of the Left is Rising to the Level of Sheer Madness #MAGA #Trump @FoxBusiness @FoxNews #Dobbs https://t.co/LTyu
WhosFibbing|t|-0.6597|0.221|0.779|0.0|RT @LouDobbs: The Ignorance of the Left is Rising to the Level of Sheer Madness #MAGA #Trump @FoxBusiness @FoxNews #Dobbs https://t.co/LTyu
NJRUA|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
BritBrat2985|realDonaldTrump|-0.6486|0.223|0.777|0.0|@realDonaldTrump @FoxNews Walking Dead is on. Watching you is the last thing I'd do Mr. Trump.
maxey_jaelen|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
carolreinoso|laurenduca|-0.5147|0.226|0.657|0.117|@laurenduca nothing gets my blood boiling more than a fellow Latino who supports Trump. WTF mi gente?!
IvanPere4|YouTube|0.0|0.0|1.0|0.0|"BREAKING: Donald Trump Just Issued Ultimatum to China! ""Do THIS or Else..."" https://t.co/l8vDwDrDT6 via @YouTube"
IvanPere4|linkis|0.0|0.0|1.0|0.0|"BREAKING: Donald Trump Just Issued Ultimatum to China! ""Do THIS or Else..."" https://t.co/l8vDwDrDT6 via @YouTube"
MarthaLivingmar|HTMLFormatNews|-0.4019|0.172|0.828|0.0|"RT @HTMLFormatNews: Clinton paid twice as much as Trump, to lose. ($1.2 billion total)https://t.co/QDpRe9BybT"
MarthaLivingmar|southjerseymechanic|-0.4019|0.172|0.828|0.0|"RT @HTMLFormatNews: Clinton paid twice as much as Trump, to lose. ($1.2 billion total)https://t.co/QDpRe9BybT"
52fairway|tribelaw|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
52fairway|twitter|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
TinaDuryea|TheDailyEdge|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
TinaDuryea|twitter|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
beyoncescurls|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
beyoncescurls||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
JeremyHimli|twitter|0.4939|0.0|0.868|0.132|"In 2008, Trump actually did work for Hillary. You know, his friend that you really thought he would  put in jail. https://t.co/HIMtponxOk"
savingfilm|sarahkendzior|0.7391|0.074|0.641|0.285|"@sarahkendzior That MSM is covering Nazis and KKK as not that bad has worked in my favor when talking to Trump supporters, weirdly."
nursiegal75|CaptainsLog2016|-0.5423|0.276|0.623|0.101|"RT @CaptainsLog2016: Dear @CanadaCan I book a 4 year stay in your country?I have no felonies, I pay taxes, and I didn't vote for Trump"
MaryTrinetti|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
CheriJacobus|twitter|0.4215|0.0|0.833|0.167|NB tweets tonight seem wisely anti-Trump even tho they don't mean them to be https://t.co/HLVsvTPUu6
Mcschweety|JoyceSt14976939|0.0|0.0|1.0|0.0|"@JoyceSt14976939 @Vis0rd0wn @KimberlyBlunk @Tim121974 @TuckerCarlson Trump can't overturn Roe V. Wade. He's president, not king."
Greg2412|JackPosobiec|-0.2168|0.161|0.719|0.12|RT @JackPosobiec: You mean like how you worked to defeat Trump's nomination? How'd that go again? https://t.co/3petpHwFvj
Greg2412|twitter|-0.2168|0.161|0.719|0.12|RT @JackPosobiec: You mean like how you worked to defeat Trump's nomination? How'd that go again? https://t.co/3petpHwFvj
KAMIAN|theslot|0.3911|0.123|0.626|0.251|"Trump Says He Doesn't Need Daily Intelligence Briefings Because He's 'You Know, Like, a Smart Person' https://t.co/hPOR4aW6gm"
PSleepyhead|JackPosobiec|0.3954|0.26|0.37|0.37|"@JackPosobiec I missed that. He did? I thought that he supported Trump. Wow, Thanks. I feel STUPID."
IntrovertRN1975|JuddLegum|-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
IntrovertRN1975||-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
Tamaraciocci|FemaleOutrage|0.0|0.0|1.0|0.0|RT @FemaleOutrage: Don't tell us that Trump wasn't coked up at the beginning of debates. Haven't heard so much sniffing since club scene in
ccarter84|StephenAtHome|-0.2714|0.165|0.712|0.124|RT @StephenAtHome: Trump has appointed a third Goldman Sachs executive to his economic team. One more and we get a free financial crisis!
lorac328|TheDailyEdge|-0.7783|0.245|0.755|0.0|RT @TheDailyEdge: Trump built his political career on the racist lie that Obama was an illegitimate President. Plot twist: he's now the ill
caroljdavy|EllenMorris1222|0.0|0.0|1.0|0.0|RT @EllenMorris1222: @JuddLegum Sucking up and covering up for Trump
KathrynGadson|alternet|0.0|0.0|1.0|0.0|5 Nightmarish Things Trump Did This Week @alternet https://t.co/kDvXIReb6m
KathrynGadson|alternet|0.0|0.0|1.0|0.0|5 Nightmarish Things Trump Did This Week @alternet https://t.co/kDvXIReb6m
librarising3|EricBoehlert|0.0|0.0|1.0|0.0|RT @EricBoehlert: Trump can't find a single senior intel official to step forward and say Russia absolutely not involved in election?
CBurtonAP|JennaFryer|0.4199|0.0|0.642|0.358|@JennaFryer that sounded Like a Trump tweet! 
cbrbwb|2ALAW|0.4048|0.0|0.786|0.214|RT @2ALAW: Isn't Christmas A Little More Special This Year? #MAGA#Trump https://t.co/o4QjFjrFEi
cbrbwb|twitter|0.4048|0.0|0.786|0.214|RT @2ALAW: Isn't Christmas A Little More Special This Year? #MAGA#Trump https://t.co/o4QjFjrFEi
A_Fellowes|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
WemittPatrick|Ramsteel007|-0.5423|0.137|0.863|0.0|RT @Ramsteel007: The CIA's SECRET plan for President TRUMP: A MUST WATCH. The CIA and MSM are enemy #2 behind Rothschild's and Soros  https
eric_walters84|MGatMES|0.4466|0.0|0.773|0.227|@MGatMES OK so what has Trump done that you say I appose?
BrownSarahM|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
TarynStanford|twitter|-0.2023|0.101|0.899|0.0|He's such a petty vindictive POS --- Trump has nailed his 'petulant 12 yr old child act.' https://t.co/PhQrrOMrx3
Read4News|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
_dsalmon|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
GettinMyWay|c0nvey|-0.0772|0.067|0.933|0.0|When Trump says he's gonna build a wall but you have a trick up your sleeve https://t.co/iFqII9pvPg by #POSITIVlBES via @c0nvey
GettinMyWay|linkis|-0.0772|0.067|0.933|0.0|When Trump says he's gonna build a wall but you have a trick up your sleeve https://t.co/iFqII9pvPg by #POSITIVlBES via @c0nvey
kaseynicolex3|TheDailyEdge|0.2263|0.087|0.791|0.123|RT @TheDailyEdge: Trump has missed 98% of his intelligence briefings. But he's always on the conference line to Moscow 5 minutes early http
eprenen|liamstack|0.0772|0.105|0.739|0.156|RT @liamstack: Now that Twitter has cracked down on the pro-Trump bots the top replies to @realDonaldTrump are mostly comedians mocking him
GarronRobert|WayneDupreeShow|0.6706|0.0|0.8|0.2|@WayneDupreeShow @Wutevuh @realDonaldTrump 2/2 irrelevant! WE NEED TO PROTECT OUR ELECTORALs! 10 4 trump are in mutiny! That is 296!
_doitfornel|GaziKodzo|0.0|0.0|1.0|0.0|RT @GaziKodzo: Trump has these white people getting they asses beat!  https://t.co/BnQtm5mkGy
_doitfornel|twitter|0.0|0.0|1.0|0.0|RT @GaziKodzo: Trump has these white people getting they asses beat!  https://t.co/BnQtm5mkGy
News4Newsman|YourAnonCentral|0.0|0.0|1.0|0.0|RT @YourAnonCentral: Democracy doesn't trump human rights. @DrHaque
SingleandSane1|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
HelenEckard|tribelaw|-0.5106|0.125|0.875|0.0|RT @tribelaw: But mounting public outrage at Trump's benefiting his family business at the expense of U.S. working men and women will do hi
MikeHighley1|Mike_Beacham|0.0|0.0|1.0|0.0|RT @Mike_Beacham: Trump says Rex Tillerson is a 'world-class player' https://t.co/0agLh4ozCk
MikeHighley1|video|0.0|0.0|1.0|0.0|RT @Mike_Beacham: Trump says Rex Tillerson is a 'world-class player' https://t.co/0agLh4ozCk
birdistheherd|260a105fb5c7455|0.2144|0.06|0.845|0.095|@260a105fb5c7455 @alfredanchor Every agency screws up and TRUMP loves to throw WMD's right in their faces but they got it RIGHT many times
AlexJHarp|katewillett|0.4767|0.0|0.86|0.14|RT @katewillett: Maybe Alec Baldwin can start reading intelligence briefings aloud on SNL to get the word to Trump somehow
AmberAufmerksam|leahmcelrath|0.0|0.0|1.0|0.0|"RT @leahmcelrath: This is a thorough compilation on @dailykos of resources regarding Putin, Dugin, Spencer, Bannon, and Trump:https://t.c"
AmberAufmerksam||0.0|0.0|1.0|0.0|"RT @leahmcelrath: This is a thorough compilation on @dailykos of resources regarding Putin, Dugin, Spencer, Bannon, and Trump:https://t.c"
dhrxsol1234|JrcheneyJohn|0.0|0.0|1.0|0.0|RT @JrcheneyJohn: The #FakeNews Media has been Neutered by Trump and they have become Irrelevant #TrumpEffect  https://t.co/8ArN8MrraK
dhrxsol1234|twitter|0.0|0.0|1.0|0.0|RT @JrcheneyJohn: The #FakeNews Media has been Neutered by Trump and they have become Irrelevant #TrumpEffect  https://t.co/8ArN8MrraK
DaveDavidmaud11|TearsInHeaven09|-0.5319|0.168|0.832|0.0|RT @TearsInHeaven09: LESSON:WHEN TRUMP TWEETS SOMETHING STUPIDHE IS TRYING TO MAKE YOU FORGETRUSSIA HACKED THE ELECTION FOR HIM
purplecait|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
MuseLotus|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
Quietness_Trust|ActionTime|-0.1531|0.144|0.743|0.114|RT @ActionTime: Please Retweet:This Must STOP-Trump's Attacks on Private Citizens on Twitter #Resist #NotMyPresident #Resistance #RT https:
prognewssource|occupydemocrats|0.25|0.067|0.817|0.115|#Breaking News: FOX Just Called Out Trump For His Pay For Play Hypocrisy To His Face https://t.co/GIr62OU6r2 by #OccupyDemocrats
mannreagan|surfermom77|-0.4215|0.128|0.872|0.0|"RT @surfermom77: The GOP bitter traitors &amp; Estab hacks, McCain &amp; Graham are joining Dems pushing the hairbrained #RussianHacking plothttps"
Sexy_Deplorable|_peripherals|-0.6229|0.185|0.815|0.0|@_peripherals maybe Trump can fix Apple too! They are ass holes and feed the liberals with their shiny toys!
rdraaf|NewYorker|0.2732|0.128|0.7|0.173|"RT @NewYorker: In the age of Trump's I love the poorly educated, Rousseau's attack on cosmopolitan lites seems prophetic. https://t.co/e"
rdraaf|twitter|0.2732|0.128|0.7|0.173|"RT @NewYorker: In the age of Trump's I love the poorly educated, Rousseau's attack on cosmopolitan lites seems prophetic. https://t.co/e"
theknottybride|EvrydayFeminism|0.4019|0.0|0.838|0.162|RT @EvrydayFeminism: We wish this didn't feel so familiar. https://t.co/bbKHO6bVeC #rapeculture #sexualassault #consent #Trump #lockerroomt
theknottybride|everydayfeminism|0.4019|0.0|0.838|0.162|RT @EvrydayFeminism: We wish this didn't feel so familiar. https://t.co/bbKHO6bVeC #rapeculture #sexualassault #consent #Trump #lockerroomt
joe_jim_regens|senrobportman|0.3182|0.0|0.881|0.119|"@senrobportman If President Elect Trump's extreme Pro Russia cabinet nominations concern you, please let Senator Portman know.  800-205-6446"
beccamarshmallo|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
beccamarshmallo||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
iggumz|FreddyLawrence1|-0.0772|0.105|0.801|0.094|"RT @FreddyLawrence1: This is spot on.It's up to @POTUS if he wants a legacy, or to have Trump finish him off being disgraced w:own party di"
gobluecoop|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
kschoon4|misscherryjones|0.0|0.0|1.0|0.0|"RT @misscherryjones: Just when I think the CIA-Russia-Trump takes can't get any hotter, along comes John Bolton with a torch."
taterpie|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
TurnTNBlue|tomtomorrow|-0.3182|0.182|0.704|0.114|"RT @tomtomorrow: Trump's  victory is as if your loved one died, and you grieve, and then they are brought back to life the next day and kil"
UcesarCesar|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
UcesarCesar|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
Run_IsHere|amjoyshow|-0.4404|0.132|0.868|0.0|"RT @amjoyshow: Scott Dworkin (@FUNDER) started #TrumpLeaks documenting hundreds of Trump's Russian ties, which the #FBI has denied or not r"
wybetter|thedailybeast|-0.7096|0.396|0.604|0.0|RT @thedailybeast: Carl Bernstein: Trump's lies worse than Nixon's:  https://t.co/wBaRkFjidX https://t.co/8lgakwPLpe
wybetter|thedailybeast|-0.7096|0.396|0.604|0.0|RT @thedailybeast: Carl Bernstein: Trump's lies worse than Nixon's:  https://t.co/wBaRkFjidX https://t.co/8lgakwPLpe
IntrovertRN1975|JuddLegum|0.128|0.0|0.897|0.103|RT @JuddLegum: 2. He's also a leading contender to be Deputy Secretary of State https://t.co/oRUPSkz7NV
IntrovertRN1975|medium|0.128|0.0|0.897|0.103|RT @JuddLegum: 2. He's also a leading contender to be Deputy Secretary of State https://t.co/oRUPSkz7NV
packergal|feliciaw5853|-0.2263|0.148|0.742|0.109|"RT @feliciaw5853: Obama trapped in presidency defining moment. Like Lincoln, unavoidable decision. Have CIA release intel on Trump. https:/"
packergal||-0.2263|0.148|0.742|0.109|"RT @feliciaw5853: Obama trapped in presidency defining moment. Like Lincoln, unavoidable decision. Have CIA release intel on Trump. https:/"
grandpooba5440|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
blueskymountain|BonhoefferLives|-0.7351|0.286|0.714|0.0|"RT @BonhoefferLives: Trump is desperately trying to distract, deny, divert, discredit the CIA, to mask his own deep complicity in nothing s"
ihaveaminutemm|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: New York Times Editorial Board demands Donald Trump go along with Russia investigation https://t.co/Fv74uavXcI via @dailynew
ihaveaminutemm|dailynewsbin|0.0|0.0|1.0|0.0|RT @starfirst: New York Times Editorial Board demands Donald Trump go along with Russia investigation https://t.co/Fv74uavXcI via @dailynew
dogmotto|Joyce_Karam|0.0|0.0|1.0|0.0|@Joyce_Karam Trump doesn't know what to say...his speechwriter on vacation.
mmsahaj|twitter|0.0|0.0|1.0|0.0|"Never wanted to talk abt Trump until now. Without evidence, we know whose side he's on. https://t.co/SWeVWf62bI"
KevinARNG11BVet|eligit|0.0|0.0|1.0|0.0|"RT @eligit: @kurteichenwald The simple fact, which has been blatantly obvious to anyone paying attention: Trump's brain cannot take in info"
ProfCAnderson|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
ProfCAnderson||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
DDianaDD|twitter|0.0|0.0|1.0|0.0| #Trump https://t.co/NJrvNrHYnv
kmh7|fightfor15|0.1027|0.165|0.652|0.183|"RT @fightfor15: (Puzder's) nomination represents the greatest assault on workers that we have seen in a generation."" https://t.co/QlQ6dEq5"
kmh7|t|0.1027|0.165|0.652|0.183|"RT @fightfor15: (Puzder's) nomination represents the greatest assault on workers that we have seen in a generation."" https://t.co/QlQ6dEq5"
Dirigo1820|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
mauree_b|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
mauree_b|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
KAMIAN|theslot|-0.0139|0.134|0.735|0.131|"Trump Says He Doesn't Need Daily Intelligence Briefings Because He's 'You Know, Like, a Sm https://t.co/lD8Tuie6oo https://t.co/kaZr1BjK50"
citizenjo|tribelaw|-0.4753|0.119|0.881|0.0|@tribelaw The thing speaks directly to Trump &amp; he still lies about it - even if it's taped! This guy is a professional conman &amp; a sociopath
nellss20|TeenVogue|-0.3612|0.185|0.815|0.0|"RT @TeenVogue: For Muslim women, a Trump presidency makes life increasingly difficult. https://t.co/9gq3zHt6c7"
nellss20|teenvogue|-0.3612|0.185|0.815|0.0|"RT @TeenVogue: For Muslim women, a Trump presidency makes life increasingly difficult. https://t.co/9gq3zHt6c7"
anthonycasey2|infowars|0.0|0.0|1.0|0.0|https://t.co/v3LTTTDisU
wtfismikeplayin|birbigs|-0.4215|0.141|0.859|0.0|RT @birbigs: Trump denies CIA report even though he doesn't read the CIA briefings...which means...wait a minute...how would he...know...th
MMaria03146111|LadyDoc4Trump|0.0|0.0|1.0|0.0|"RT @LadyDoc4Trump: Our ""president"" says NOTHING, NADA, ZERO about #Christian genocide by his Muslim brothers.#Trump speaks #Truth on it."
Jennuendoh|OhNoSheTwitnt|-0.7003|0.254|0.746|0.0|"RT @OhNoSheTwitnt: A game called ""Actual Trump Tweet or Parody Account?"" and you lose whether you guess right or wrong."
honorverity|Gundlefinger16|0.6369|0.101|0.57|0.329|RT @Gundlefinger16: @Khanoisseur She would be a great president. Trump interrupts to prevent the truth from coming out.
RachelK1967|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Ltr from Hon Elijah Cummings asking Chaffetz to Investigate Trump biz conflicts#cnn #msnbc #AMJoy #cnnsotu #this
sf49ersfan5249|LouDobbs|-0.6597|0.221|0.779|0.0|RT @LouDobbs: The Ignorance of the Left is Rising to the Level of Sheer Madness #MAGA #Trump @FoxBusiness @FoxNews #Dobbs https://t.co/LTyu
sf49ersfan5249|t|-0.6597|0.221|0.779|0.0|RT @LouDobbs: The Ignorance of the Left is Rising to the Level of Sheer Madness #MAGA #Trump @FoxBusiness @FoxNews #Dobbs https://t.co/LTyu
AdvocatAmy1|howiewolf|0.0|0.0|1.0|0.0|RT @howiewolf: Emails found on Anthony Weiner's computer? Tell the world. Russians trying to elect Donald Trump? Sweep it under the rug.
jyester55|LawyerRogelio|-0.7034|0.277|0.639|0.084|RT @LawyerRogelio: NYC DISLIKES TRUMPS Supposedly tolerant NYC is making the Trump kids lives horrible | New York Post https://t.co/rP5g
jyester55|t|-0.7034|0.277|0.639|0.084|RT @LawyerRogelio: NYC DISLIKES TRUMPS Supposedly tolerant NYC is making the Trump kids lives horrible | New York Post https://t.co/rP5g
statefarm2005|MSNBC|0.2057|0.0|0.932|0.068|@MSNBC The media is not biased against Trump. All they are doing is reporting on what he does. Same with Clinton. They report what she does.
gbeckyhudson|bourgeoisalien|-0.6656|0.214|0.786|0.0|"RT @bourgeoisalien: Trump said he doesn't need intelligence briefings bc he's 'smart' yet watches news he hates daily. Um, 'smart' isn't yo"
chrissmax|facebook|0.9022|0.0|0.59|0.41|Trump loves Russia. Russia loves Trump. So let's make everyone happy and have Trump be President of Russia. https://t.co/DMYDauuejJ
simi_kc88|USARedOrchestra|0.0|0.0|1.0|0.0|"RT @USARedOrchestra: CT Rep. Jim Himes call Trump ""completely unhinged"" and calls for the electoral college to do what it was designed for."
Hope_NoelB|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
PatPatojson|Corporatocrazy|-0.8316|0.328|0.672|0.0|"RT @Corporatocrazy: Two things CIA could be doing now:A. Kill ISIS, orB. Spread fake news to delegitimize Trumphttps://t.co/RzTTRpgvp8"
BigBobGardner|nytimes|0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
BigBobGardner||0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
AmesCG|JohnFPfaff|-0.0516|0.095|0.905|0.0|"RT @JohnFPfaff: So if each daily briefing says ""Russians are ten miles closer to Warsaw than yesterday,"" how long after Warsaw falls will T"
DebbieW36246900|TeeTweetsHere|-0.802|0.324|0.676|0.0|"RT @TeeTweetsHere: In Response To Hate Crime Spike, Muslim NYPD Officers Ask For Meeting With Trump https://t.co/2WamQ9JOaV"
DebbieW36246900|huffingtonpost|-0.802|0.324|0.676|0.0|"RT @TeeTweetsHere: In Response To Hate Crime Spike, Muslim NYPD Officers Ask For Meeting With Trump https://t.co/2WamQ9JOaV"
barney_cannon|TeaPainUSA|0.128|0.092|0.797|0.112|"RT @TeaPainUSA: Trump claims the CIA said Saddam had WMDs.  Ironically, he's thinkin' of the last President that lost the popular vote."
SscottSsmith84|DrEstella|0.0|0.0|1.0|0.0|"RT @DrEstella: Senator #HarryRead asks CIA to lie to @realDonaldTrump ""Give Trump ""Fake"" INTEL BRIEFINGS!""  #SundayMorning #WeareTrump #Tru"
Hot_Techie_News|hottechienews|-0.4019|0.267|0.593|0.141|Donald Trump Clarifies His Plans for Destroying theEnvironment https://t.co/KBW3GuZjZS https://t.co/hrdMptC7Tx
PaulJon54388869|swin24|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
PaulJon54388869|thedailybeast|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
bristow72|kellwoohoo|0.0|0.0|1.0|0.0|RT @kellwoohoo: Translation: Trump will appoint people who'll look the other way &amp; let Russia get away with anything &amp; everything. https://
bristow72||0.0|0.0|1.0|0.0|RT @kellwoohoo: Translation: Trump will appoint people who'll look the other way &amp; let Russia get away with anything &amp; everything. https://
barSwilson|linkis|0.0|0.0|1.0|0.0|"Drumpf: I'd 'love' to have Ivanka, Jared Kushner 'involved' https://t.co/gxgZiM1uqW"
CraigSymons|seanmdav|0.4728|0.044|0.836|0.12|"RT @seanmdav: A stray thought: if media didn't want Trump in the WH, perhaps they shouldn't have showered him w/ $2 billion in free GOP pri"
Twinmommie09|change|-0.296|0.196|0.804|0.0|Petition update - You Can Stop Trump on December 19 https://t.co/G9ukRd5tLQ
TheDailyDigest|newfoundland|0.0|0.0|1.0|0.0|"Trump calls Russian election influence report ""ridiculous"" https://t.co/9TSQyV2wEL"
Celebrilizer|celebs|0.0|0.0|1.0|0.0|Trump: I'd 'Love' to Have #IvankaInvolved in Administration #JaredKushner #DonaldTrump https://t.co/J70y31CrWW https://t.co/jgYTgMDSO8
maegabby49|JuddLegum|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
maegabby49|medium|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
Maxzen2004|Vote_American|0.0|0.0|1.0|0.0|"RT @Vote_American: @AmyMek @826Maureen @realDonaldTrump Today, Trump Made a Chump Out of Obama Today! By Attending the Army/Navy Game! http"
TRUMPIS4US|JackPosobiec|-0.2168|0.161|0.719|0.12|RT @JackPosobiec: You mean like how you worked to defeat Trump's nomination? How'd that go again? https://t.co/3petpHwFvj
TRUMPIS4US|twitter|-0.2168|0.161|0.719|0.12|RT @JackPosobiec: You mean like how you worked to defeat Trump's nomination? How'd that go again? https://t.co/3petpHwFvj
steveg1425|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
iamjoemeyer|BettyBowers|0.0|0.0|1.0|0.0|"RT @BettyBowers: If I write something about Trump &amp; you respond by digging up a worn-out meme about Clinton or Obama, youre saying, I can"
joh53293471|MissPride2u|0.5423|0.088|0.683|0.229|"RT @MissPride2u: Dear Electoral College, The fact that Donald Trump refused intelligence briefings should give you food for thought. Vote @"
burberryant|jring383|0.3182|0.0|0.874|0.126|RT @jring383: @dshanesmith @billmaher since when does wanting a fresh face for a progressive agenda synonymous with embracing Trump?
IntrovertRN1975|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
IntrovertRN1975|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
Paidsubscriber|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
WilliamSnowHume|yugvaniworld|-0.5106|0.155|0.845|0.0|@yugvaniworld And TRUMP rejected the CIA long before the election.  Here's why he was right to do that:  https://t.co/afU0DjTiHG
WilliamSnowHume|cnn|-0.5106|0.155|0.845|0.0|@yugvaniworld And TRUMP rejected the CIA long before the election.  Here's why he was right to do that:  https://t.co/afU0DjTiHG
Sheilas11|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
1775reaper|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: Trump: 'Nobody really knows' if #ClimateChange is real. Um... Apart from every scientist who works on the subject?! Idi
sudnapo|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
stanthemanchan|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
Cantuono|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
gabbysherrill|realDonaldTrump|0.8478|0.0|0.595|0.405|"@realDonaldTrump @NBCNightlyNews @CNN Praying for you daily, President Trump. Please stay focused. We are on your side. Thank you!"
Panther_NoTiger|NAVolatPropriis|0.1027|0.159|0.619|0.221|"RT @NAVolatPropriis: I just feel like in every other space, a person acting like Trump would have been fired."
mapnotes|jerryaldeeni|0.0|0.0|1.0|0.0|RT @jerryaldeeni: https://t.co/CxzMzmql8z
mapnotes|nytimes|0.0|0.0|1.0|0.0|RT @jerryaldeeni: https://t.co/CxzMzmql8z
danfelix82|Lglwry|-0.6114|0.182|0.818|0.0|"@Lglwry @HeideggerFan @justinhendrix hey dummy, not one agency has implied Trump was involved at all.  Wishful thinking yet pathetic!"
writeshawn|glennspizza|-0.1027|0.167|0.833|0.0|"RT @glennspizza: ""maggie for president"" trump is shook"
RhapsodysBIues|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
springerthings|misscherryjones|0.0|0.0|1.0|0.0|"RT @misscherryjones: Just when I think the CIA-Russia-Trump takes can't get any hotter, along comes John Bolton with a torch."
carnifexia|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
whinknee|Salon|-0.743|0.283|0.717|0.0|RT @Salon: 3 people on Trump's team have been accused of physical or sexual violence against women https://t.co/tsY1Pb5PSU https://t.co/9iF
whinknee|salon|-0.743|0.283|0.717|0.0|RT @Salon: 3 people on Trump's team have been accused of physical or sexual violence against women https://t.co/tsY1Pb5PSU https://t.co/9iF
PercyChekov|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
PercyChekov|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
MikaelaSkyeSays|kurteichenwald|-0.5423|0.176|0.824|0.0|"RT @kurteichenwald: Fox/Cheney went nuts when found out Obama got intel briefings in writing, rather than read to him. But Trump no briefin"
Rene2608|twitter|-0.6571|0.522|0.478|0.0|That's right!!! Fuck Trump  https://t.co/bZn8OotP7k
Betsyg6Gervasi|USARedOrchestra|0.0|0.0|1.0|0.0|"RT @USARedOrchestra: CT Rep. Jim Himes call Trump ""completely unhinged"" and calls for the electoral college to do what it was designed for."
MissUSA56|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
JonSteege|JuddLegum|-0.4939|0.167|0.833|0.0|RT @JuddLegum: Donald Trump confirms he will violate the Constitution on his first day in office https://t.co/CEW1XUMbeV
JonSteege|medium|-0.4939|0.167|0.833|0.0|RT @JuddLegum: Donald Trump confirms he will violate the Constitution on his first day in office https://t.co/CEW1XUMbeV
deymartin|twitter|-0.5267|0.207|0.793|0.0|Electors must do the right thing. Donald Trump is a danger to our republic. https://t.co/VDDOnCZSFs
Jrjaja1|DENVERSMKC|0.0|0.0|1.0|0.0|@DENVERSMKC @JoyAnnReid Hey this is just d beginning. Trump isn't going 2bsatisfied w a few millions. We r talking about multi Billions NOW
Neethz426|AlecBaldwin|0.8065|0.0|0.658|0.342|Best Guest Performer in a Comedy Series - @AlecBaldwin for his Trump impersonation on @nbcsnl !! #CriticsChoice https://t.co/fMEnVROm68
Neethz426|twitter|0.8065|0.0|0.658|0.342|Best Guest Performer in a Comedy Series - @AlecBaldwin for his Trump impersonation on @nbcsnl !! #CriticsChoice https://t.co/fMEnVROm68
carolyn_pearl|SenSanders|0.4767|0.08|0.691|0.229|"RT @SenSanders: I challenge Mr. Trump to tell the American people he'll keep his promises and veto cuts to Social Security, Medicare and Me"
OnceUpo00786525|npr|0.0|0.0|1.0|0.0|via @npr: CIA Concludes Russian Interference Aimed To Elect Trump https://t.co/tg3MUcxSoc
OnceUpo00786525|npr|0.0|0.0|1.0|0.0|via @npr: CIA Concludes Russian Interference Aimed To Elect Trump https://t.co/tg3MUcxSoc
bluebonnetbunny|DMansini|0.4926|0.0|0.814|0.186|RT @DMansini: Trump Jr. Held Secret Talks With Russia Supporters https://t.co/AsGZU1Ov1u via @thedailybeastENOUGH! #InvestigateTrumpNOW @T
bluebonnetbunny|thedailybeast|0.4926|0.0|0.814|0.186|RT @DMansini: Trump Jr. Held Secret Talks With Russia Supporters https://t.co/AsGZU1Ov1u via @thedailybeastENOUGH! #InvestigateTrumpNOW @T
Tull007|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
Tull007|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
2figures2|V_of_Europe|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
2figures2|thegatewaypundit|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
themanamedan|twitter|0.0|0.0|1.0|0.0|How long until it's trump https://t.co/AtO2Wof8xJ
JoinerMari|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS: GOP on hill ""prepping for President Pence""-Trump investigation begins-More soon#cnn #msnbc #AMJoy #cnnsotu #this"
Regency_Reader|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
AlpalCarla|SocialPowerOne1|0.3182|0.111|0.702|0.187|RT @SocialPowerOne1: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests https://t.co/Eghd6ic7s8
AlpalCarla|politicususa|0.3182|0.111|0.702|0.187|RT @SocialPowerOne1: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests https://t.co/Eghd6ic7s8
TNChick67|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Uncovered-Before Donald Trump Made A Deal With Carrier, He Sued It@JoyAnnReid #obama #msnbc #cnn #dnc https://t.c"
TNChick67||0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Uncovered-Before Donald Trump Made A Deal With Carrier, He Sued It@JoyAnnReid #obama #msnbc #cnn #dnc https://t.c"
ToWoods|mariabustillos|-0.5423|0.242|0.641|0.117|RT @mariabustillos: Some backstory on bad novelist and gigantic idiot Ayn Rand (so beloved of Trump cabinet) that I wrote @Awl https://t.co
ToWoods|t|-0.5423|0.242|0.641|0.117|RT @mariabustillos: Some backstory on bad novelist and gigantic idiot Ayn Rand (so beloved of Trump cabinet) that I wrote @Awl https://t.co
valeriobrl|NYCMayor|0.0|0.0|1.0|0.0|@NYCMayor   Finds His Mojo as the Anti-Trump https://t.co/TLzqMRziVL
valeriobrl|politico|0.0|0.0|1.0|0.0|@NYCMayor   Finds His Mojo as the Anti-Trump https://t.co/TLzqMRziVL
mausiepup|MarkHarrisNYC|-0.8555|0.331|0.669|0.0|RT @MarkHarrisNYC: Those briefings scare Trump--they're full of info he doesn't know and can't hold onto. And being scared angers him.  htt
caroljdavy|JuddLegum|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
caroljdavy|medium|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
Gjizzle55|yashar|0.0|0.0|1.0|0.0|"RT @yashar: WATCH: Trump's expected nominee for Deputy Secretary of State, John Bolton, trashing the UN and wading in a pool of nationalism"
DaveJRosas|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
DaveJRosas|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
CountryLiberal|pattonoswalt|0.4939|0.076|0.763|0.16|RT @pattonoswalt: Donald Trump has made me re-consider my love of Rodney Dangerfield's character in CADDYSHACK and for that alone he should
winkiechance|slone|0.8176|0.0|0.691|0.309|RT @slone: #GOPe House &amp; Senate better understand that @realDonaldTrump supporters do NOT support them &amp; their BS GLOBALIST agenda. We supp
JohnPietaro|moveon|0.3818|0.0|0.852|0.148|Independent Caucus NY Senate Democrats Must Unite to Protect NY State from Donald Trump https://t.co/8oyGrkfEfk @moveon
JohnPietaro|petitions|0.3818|0.0|0.852|0.148|Independent Caucus NY Senate Democrats Must Unite to Protect NY State from Donald Trump https://t.co/8oyGrkfEfk @moveon
Lucy59jarvis|immigrant4trump|0.6588|0.0|0.82|0.18|RT @immigrant4trump: Video: Trump is going to Make America Great Again Regardless of the Color of your Skin! #Maga #Trump https://t.co/3aDj
Lucy59jarvis|t|0.6588|0.0|0.82|0.18|RT @immigrant4trump: Video: Trump is going to Make America Great Again Regardless of the Color of your Skin! #Maga #Trump https://t.co/3aDj
TonyHui99|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
TonyHui99|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
blingdomepiece|jnpaquet|0.34|0.0|0.897|0.103|RT @jnpaquet: Norwegian cartoonist Christian Bloom is creator of this cartoon of #Trump that has recently been shared on Twitter before cen
dr_ashok_m|joshob1987|0.25|0.172|0.594|0.234|RT @joshob1987: Because they have to present it like they are definitely sure Russia rigged it for Trump &amp; they must be attacked immediatel
metroadlib|DavidCornDC|0.0|0.0|1.0|0.0|RT @DavidCornDC: Why Donald Trump appointing John Bolton to any post is crazy...even for Trump: https://t.co/KjbZP4B4Z3
metroadlib|m|0.0|0.0|1.0|0.0|RT @DavidCornDC: Why Donald Trump appointing John Bolton to any post is crazy...even for Trump: https://t.co/KjbZP4B4Z3
Myop1357|amjoyshow|-0.5267|0.139|0.861|0.0|RT @amjoyshow: .@TRIBELAW says due to emoluments clause: The Constitution is going to be violated the moment #Trump takes the oath. RETWEET
ToddDomke|BrendanNyhan|0.0|0.0|1.0|0.0|RT @BrendanNyhan: Reminder: Trump has not disclosed finances that could reveal Russian ties &amp; could be enriched by them via businesses now
thebobbyb|MrDane1982|-0.2808|0.172|0.71|0.118|"RT @MrDane1982: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/osh9DydG9E via @Bipartisan"
thebobbyb|bipartisanreport|-0.2808|0.172|0.71|0.118|"RT @MrDane1982: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/osh9DydG9E via @Bipartisan"
SandraDighton1|infidel_murdoc|0.6166|0.0|0.817|0.183|@infidel_murdoc YOU TRUST TRUMP RE BUY AMERICA HIRE AMERICA WHEN HE JUST APPLIED FOR WORK VISAS FOR MIR LAGO
FunnyFaceKing|MartinShovel|0.3182|0.0|0.796|0.204|RT @MartinShovel: My cartoon - Truth vs Post-Truth#Brexit #Trump #r4Today  https://t.co/uPeaokus2z
FunnyFaceKing|twitter|0.3182|0.0|0.796|0.204|RT @MartinShovel: My cartoon - Truth vs Post-Truth#Brexit #Trump #r4Today  https://t.co/uPeaokus2z
wildwonderweb|SeanMcElwee|0.0|0.0|1.0|0.0|RT @SeanMcElwee: *Trump appoints six of his biggest donors to high-ranking cabinet positions*New York Times: https://t.co/6nDnnrBh85
wildwonderweb|twitter|0.0|0.0|1.0|0.0|RT @SeanMcElwee: *Trump appoints six of his biggest donors to high-ranking cabinet positions*New York Times: https://t.co/6nDnnrBh85
shiphitsthefan|SarcasticRover|0.0|0.0|1.0|0.0|RT @SarcasticRover: ALL THE F--KING SCIENTISTS KNOW. https://t.co/NMqukcqfme
shiphitsthefan|washingtonpost|0.0|0.0|1.0|0.0|RT @SarcasticRover: ALL THE F--KING SCIENTISTS KNOW. https://t.co/NMqukcqfme
Smize21|ButchJocson|0.7249|0.0|0.789|0.211|"RT @ButchJocson: 62+million Americans voted for Donald J Trump, influenced &amp; behooved by a very simple common sense love for the USA!!!"
magpie51pa|ClimateReality|0.5994|0.0|0.776|0.224|"RT @ClimateReality: #DYK? In some parts of the United States, wind energy is the cheapest electricity source available https://t.co/OdhDVYc"
magpie51pa|t|0.5994|0.0|0.776|0.224|"RT @ClimateReality: #DYK? In some parts of the United States, wind energy is the cheapest electricity source available https://t.co/OdhDVYc"
FMAlchemist|RawStory|-0.34|0.124|0.876|0.0|"RT @RawStory: Foxs Judge Jeanine has bonkers rant: If you investigate Russian 2016 hacking, youre against America https://t.co/iTENvK7MKC"
FMAlchemist|rawstory|-0.34|0.124|0.876|0.0|"RT @RawStory: Foxs Judge Jeanine has bonkers rant: If you investigate Russian 2016 hacking, youre against America https://t.co/iTENvK7MKC"
Weshauk|WSJ|-0.4767|0.341|0.659|0.0|@WSJ @johndmckinnon Trump means for himself. Shame
afinndorian|realDonaldTrump|0.3595|0.0|0.858|0.142|"@realDonaldTrump President Trump will restore Manhood in this Country, leading by example.Accountability is going to return!"
TheResi12243329|CeeLeeMusic|0.0|0.0|1.0|0.0|RT @CeeLeeMusic: People keep saying Trump picked #Tillerson for SOS.No. Let's be clear.Vladimir Putin picked Tillerson.#RussianHacker
lonegamer78|pattonoswalt|-0.2732|0.196|0.675|0.129|RT @pattonoswalt: Well shithouse mouse. @TeenVogue nails the frightening absurdity of Trump... https://t.co/d8mKBjmGDL
lonegamer78|twitter|-0.2732|0.196|0.675|0.129|RT @pattonoswalt: Well shithouse mouse. @TeenVogue nails the frightening absurdity of Trump... https://t.co/d8mKBjmGDL
ElaineCarlisl1|ElaineCarlisl1|0.6688|0.0|0.766|0.234|RT @ElaineCarlisl1: Attention Trump fans! Donald Trump is giving you a lesson on how to style your hair like him! https://t.co/CO87iJPUuu
ElaineCarlisl1|twitter|0.6688|0.0|0.766|0.234|RT @ElaineCarlisl1: Attention Trump fans! Donald Trump is giving you a lesson on how to style your hair like him! https://t.co/CO87iJPUuu
AmyZanrosso|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
biotrooferredux|DarthPutinKGB|0.0|0.0|1.0|0.0|"RT @DarthPutinKGB: By the time you've figured out what we did to get Trump elected, we'll have overthrown Merkel."
EnriqueM77|Cernovich|0.103|0.079|0.787|0.134|"RT @Cernovich: Trump is not a perfect man, flawed to be sure like everyone else, but compared to Clintons (either of them), he's a saint."
jmingerson725|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
wmikenelson|ejenk|0.7906|0.0|0.696|0.304|RT @ejenk: I saw a video of Russians cheering on the rooftops in New Jersey when Trump won the election.
Donaldson2016|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
Donaldson2016|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
dnparkerson|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
dnparkerson||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
mauree_b|JuddLegum|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
mauree_b|medium|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
caroljdavy|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
caroljdavy|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
zacnba|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
am_goed|SarahPalinUSA|-0.0422|0.118|0.77|0.112|RT @SarahPalinUSA: Russia's getting out of hand? So says the defeated. Not to worry... remember I can keep an eye on them from here. https:
pamelaval|Truth2Power2016|0.0|0.0|1.0|0.0|@Truth2Power2016 @ArmyVet64 @MelissaJPeltier @MagicManArthur Trump colluded says the agenda-laden MSM.  Hilary collided selling 20% uranium
Pu55yGalore|TeaPainUSA|0.34|0.0|0.893|0.107|"RT @TeaPainUSA: Trump says security briefings say the same thing every day: ""Putin has compromised multiple positions at the highest level"
pjcags|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
pjcags||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
kp_ppkp2013|TIME|0.0|0.0|1.0|0.0|RT @TIME: Meet the voters who helped put Donald Trump in the White House #TIMEPOY https://t.co/fW1FwQefng
kp_ppkp2013|time|0.0|0.0|1.0|0.0|RT @TIME: Meet the voters who helped put Donald Trump in the White House #TIMEPOY https://t.co/fW1FwQefng
BerneStober|AP4LP|0.3244|0.0|0.885|0.115|"RT @AP4LP: Liberal Logic: ""You dont need assault rifles. Govt wont turn tyrannical but Trump is the next Hitler!"""
acidddsaint|acidddsaint|-0.3182|0.119|0.881|0.0|RT @acidddsaint: do you guys think that if trump lost a little bit of weight...maybe his neck will emerge?
nytrb|nytimes|0.0|0.0|1.0|0.0|Trump Suggests Using Bedrock China Policy as Bargaining Chip - New York Times https://t.co/jyMdvhzFYj
Tull007|JuddLegum|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
Tull007|medium|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
TheKidRosenbaum|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
TheKidRosenbaum|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
carolinelv|thehill|0.0|0.0|1.0|0.0|RT @thehill: Christie turned down several positions in Trump administration: reporthttps://t.co/Ff4dxZ0zkz https://t.co/LVefpPfmiC
carolinelv|twitter|0.0|0.0|1.0|0.0|RT @thehill: Christie turned down several positions in Trump administration: reporthttps://t.co/Ff4dxZ0zkz https://t.co/LVefpPfmiC
verarocks|ryanlips|0.0|0.0|1.0|0.0|RT @ryanlips: Reboot of Mystery Science Theater 3000 but the robots are Donald Trump and the movies are the news.
tin_10001|business|-0.34|0.167|0.833|0.0|RT @business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/6l8izhUs9D https://t.co/0drSTTUrnr
tin_10001|bloomberg|-0.34|0.167|0.833|0.0|RT @business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/6l8izhUs9D https://t.co/0drSTTUrnr
Gjizzle55|nytimes|0.0|0.0|1.0|0.0|"RT @nytimes: Boeing Seeks to Sell Planes to Iran, and the Deal to Trump https://t.co/VsnlIkl4Ss"
Gjizzle55|nytimes|0.0|0.0|1.0|0.0|"RT @nytimes: Boeing Seeks to Sell Planes to Iran, and the Deal to Trump https://t.co/VsnlIkl4Ss"
chicashawna|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
brady_aol|richardharris69|0.1027|0.118|0.746|0.136|RT @richardharris69: BREAKING NEWS:  an investigation has found that Trump skips intelligence briefings because he has a problem with the w
tomphillipsin|JohnDelury|-0.7469|0.189|0.811|0.0|"RT @JohnDelury: Not to be alarmist, but when I asked what Beijing will do if Trump persists w Two China Policy, the answer was war https://"
tomphillipsin||-0.7469|0.189|0.811|0.0|"RT @JohnDelury: Not to be alarmist, but when I asked what Beijing will do if Trump persists w Two China Policy, the answer was war https://"
petrified_syrup|TheDailyEdge|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
petrified_syrup|twitter|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
JulieMcGill11|asamjulian|-0.1027|0.055|0.945|0.0|"RT @asamjulian: Chris Wallace says Trump is ""almost more the president than the president is"" and that we pay more attention to him than Ob"
joehoevah|micahcohen|-0.8519|0.377|0.623|0.0|"RT @micahcohen: How much harm is done, in media and government, from the fear of being accused of bias? https://t.co/zkcp9an5Oi https://t.c"
joehoevah|nytimes|-0.8519|0.377|0.623|0.0|"RT @micahcohen: How much harm is done, in media and government, from the fear of being accused of bias? https://t.co/zkcp9an5Oi https://t.c"
blahblahellis|twitter|0.0|0.0|1.0|0.0|"They put a bit of coal in Kirk Douglass's fist and said: ""Trump"". https://t.co/Yc1UqmeDoA"
WePeople2016|thehill|-0.4404|0.195|0.805|0.0|"RT @thehill: SNL fires back at Trump criticism: We know ""he's watching""https://t.co/3Y5IM7U35z https://t.co/KCW8AZ8y9r"
WePeople2016|thehill|-0.4404|0.195|0.805|0.0|"RT @thehill: SNL fires back at Trump criticism: We know ""he's watching""https://t.co/3Y5IM7U35z https://t.co/KCW8AZ8y9r"
NTrexit|Change|-0.4404|0.255|0.607|0.138|US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/XXcabkIMcP via @Change
NTrexit|change|-0.4404|0.255|0.607|0.138|US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/XXcabkIMcP via @Change
JaneGummyof3|HamiltonElector|0.2298|0.123|0.757|0.12|"RT @HamiltonElector: Mr. Trump you are hardly a genius, no matter what Comrade Putin says.  We are smarter than you. We are #hamiltonelecto"
AugustEve2012|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
PaulJon54388869|swin24|-0.0572|0.055|0.945|0.0|"RT @swin24: Today, Trump says he doesnt want anyone hacking the U.S.In July, he called on Russia to hack the U.S. govt.https://t.co/"
pamplemoussee76|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
smokestacklite|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Ltr from Hon Elijah Cummings asking Chaffetz to Investigate Trump biz conflicts#cnn #msnbc #AMJoy #cnnsotu #this
grandpooba5440|KeithOlbermann|-0.4588|0.13|0.87|0.0|"RT @KeithOlbermann: CIA says Russia intervened to elect Trump. Trump sides with Russia, mocks CIA. From 11/1: The Trumpchurian Candidate ht"
fool4thetruth|twitter|-0.8225|0.336|0.664|0.0|Russia wanted Trump to win?Maybe they did to avert Nuclear War that Hillary threatened them with her WHOLE CAMPAIGN https://t.co/aZNQHEWQUw
RedRose3b|RadioFreeTom|0.4767|0.0|0.876|0.124|"RT @RadioFreeTom: If HRC chose a SecState who ran an oil giant and got a medal from Putin, the GOPers defending Trump would re-convene the"
Lina_J_Al|anders_aslund|-0.8834|0.424|0.576|0.0|"RT @anders_aslund: @SenJohnMcCain hitting hard: ""Vladimir Putin is a thug and a murderer and a killer and a KGB agent. https://t.co/Itkjg4"
Lina_J_Al|t|-0.8834|0.424|0.576|0.0|"RT @anders_aslund: @SenJohnMcCain hitting hard: ""Vladimir Putin is a thug and a murderer and a killer and a KGB agent. https://t.co/Itkjg4"
clark7950|SpecialKMB1969|0.4019|0.0|0.847|0.153|RT @SpecialKMB1969: Just picked up the November's @Newsweek Special Commemorative EditionPRESIDENT TRUMP #Newsweek DJT's Historic Journey
jmhodges|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
jmhodges|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
wtf_imtooold|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
Bay_St_Wiseguy|CarmineZozzora|-0.6486|0.218|0.782|0.0|"RT @CarmineZozzora: Everything we've witnessed the last 19 months, and including today's Russian fake news narrative, has been coup to stop"
trishmaximum|blockchainhelpr|-0.296|0.128|0.872|0.0|RT @blockchainhelpr: Are You Worried About Trump? Then Start Your Own Country #donaldtrump #blockchain https://t.co/uVxBSw7GGP https://t.co
trishmaximum|blockgeeks|-0.296|0.128|0.872|0.0|RT @blockchainhelpr: Are You Worried About Trump? Then Start Your Own Country #donaldtrump #blockchain https://t.co/uVxBSw7GGP https://t.co
AnitaStubbs|HamiltonElector|-0.296|0.099|0.901|0.0|RT @HamiltonElector: We've crossed the threshold. There is no going back. Trump must never become POTUS. RT to let #hamiltonelectors know y
Bayathread|feministing|0.5859|0.0|0.703|0.297|@feministing follow @RachelleHodgs for brilliant graphing of Trump word salads.
richiebel|Will_Bunch|-0.7149|0.239|0.761|0.0|"RT @Will_Bunch: Worse than Watergate? Russia hacking is massive cloud over Trump presidency, and America. What caused this big mess? https:"
Ivy_B|Will_Bunch|-0.7149|0.239|0.761|0.0|"RT @Will_Bunch: Worse than Watergate? Russia hacking is massive cloud over Trump presidency, and America. What caused this big mess? https:"
RockyinTX|rjoseph7777|-0.7096|0.396|0.604|0.0|RT @rjoseph7777: Bernstein: Trumps Lies Worse Than Nixons  https://t.co/kup1gmrE13 #RussiaHacking #Unfit
RockyinTX|thedailybeast|-0.7096|0.396|0.604|0.0|RT @rjoseph7777: Bernstein: Trumps Lies Worse Than Nixons  https://t.co/kup1gmrE13 #RussiaHacking #Unfit
princessmom122|matthewjdowd|0.0|0.0|1.0|0.0|"RT @matthewjdowd: So Trump knows more about business than Wall Street Journal, more about military than Generals, and more about intelligen"
jewbaby57|Democrat_4Trump|-0.516|0.305|0.461|0.234|RT @Democrat_4Trump: Teacher Calls Trump Win TERRORISM: Caught On Hidden Camera Calling Trump Win An 'Act Of Terrorism' https://t.co/QYoqa9
jewbaby57|t|-0.516|0.305|0.461|0.234|RT @Democrat_4Trump: Teacher Calls Trump Win TERRORISM: Caught On Hidden Camera Calling Trump Win An 'Act Of Terrorism' https://t.co/QYoqa9
SalatapNagol15|MattWalshBlog|0.0|0.0|1.0|0.0|RT @MattWalshBlog: The fact is this: Russia didn't elect Donald Trump. The American people did.
AuerbachKeller|adamjohnsonNYC|0.0516|0.132|0.726|0.141|RT @adamjohnsonNYC: during the primaries it was real news--not fake news--that gave Trump $1.8 billion in free media https://t.co/dSuiSWRjj
AuerbachKeller|t|0.0516|0.132|0.726|0.141|RT @adamjohnsonNYC: during the primaries it was real news--not fake news--that gave Trump $1.8 billion in free media https://t.co/dSuiSWRjj
RenoSteph|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
BlakeGordon17|andieiamwhoiam|0.5267|0.065|0.75|0.185|"RT @andieiamwhoiam: Sorry Lefties, Russians, recounts, aliens (the extraterrestrial kind)...you will never get a new election.  Trump won."
Sugalean|davepell|-0.7713|0.22|0.745|0.036|"RT @davepell: No matter what the Russians did, the most devastating story of 2016 is that Americans saw Trump for what he is and voted for"
Fernasteady|Evan_McMullin|-0.1027|0.129|0.759|0.112|"RT @Evan_McMullin: Trump encouraged Russian subversion of our democracy then denied its occurrence despite CIA evidence, while preparing to"
lonegamer78|pattonoswalt|-0.5719|0.209|0.791|0.0|RT @pattonoswalt: And then @TeenVogue illustrates the horror of Trump's America on the ground... https://t.co/2ZLaIuA15y
lonegamer78|twitter|-0.5719|0.209|0.791|0.0|RT @pattonoswalt: And then @TeenVogue illustrates the horror of Trump's America on the ground... https://t.co/2ZLaIuA15y
Who_R_U82|Lilliana1017|-0.5719|0.222|0.778|0.0|RT @Lilliana1017: Someone keeps photoshopping Trump's face on the Queen and it's terrifying https://t.co/4wsO3aLUVg
Who_R_U82|yahoo|-0.5719|0.222|0.778|0.0|RT @Lilliana1017: Someone keeps photoshopping Trump's face on the Queen and it's terrifying https://t.co/4wsO3aLUVg
sud_vijay|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
oursisthehour|stanleyrogouski|-0.1027|0.174|0.714|0.112|RT @stanleyrogouski: Do the Democrats actually believe they're going to stop Trump by accusing him of being a Russian asset?
RamsenRasho|ImpeachPOTUS|0.6249|0.0|0.745|0.255|@ImpeachPOTUS @Jennifer4130 shut your mouth and watch trump make America great again bimbo.
FededelCorro|vickytedije|0.4588|0.0|0.842|0.158|"@vickytedije viendo los People Choice awards entends que haya ganado Trump y Macri, la gente vota cualquier cosa."
colbert_ed|davidfrum|0.7351|0.0|0.754|0.246|"RT @davidfrum: US intelligence community: Russia acted to install Trump. 18 months from now, there wont be a US intelligence community wor"
mminajohnson|andylassner|0.0431|0.123|0.713|0.163|RT @andylassner: Do NOT use this photo of Donald Trump. He does NOT like it. He told reporters he HATES it. Please RETWEET. https://t.c
mminajohnson||0.0431|0.123|0.713|0.163|RT @andylassner: Do NOT use this photo of Donald Trump. He does NOT like it. He told reporters he HATES it. Please RETWEET. https://t.c
lsuagain|PSheritaakkloh|-0.6199|0.238|0.762|0.0|"@PSheritaakkloh @Ckzoote If you hate Trump, why are you following his tweets? Troll much?"
DomAcconcia|politico|0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
DomAcconcia||0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
SusanIverach|WeNeedTrump|0.0|0.0|1.0|0.0|RT @WeNeedTrump: BOOM: Look at the LOCKER ROOM dedication they gave Trump at the Army/Navy game!https://t.co/dc0HEwjZ0L
SusanIverach|ilovemyfreedom|0.0|0.0|1.0|0.0|RT @WeNeedTrump: BOOM: Look at the LOCKER ROOM dedication they gave Trump at the Army/Navy game!https://t.co/dc0HEwjZ0L
rbean14620|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
rbean14620|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
DAILYBLUEblog|sarahkendzior|-0.296|0.109|0.891|0.0|"RT @sarahkendzior: In the ever-evolving shakedown, Trump is peddling an ""Inaugural Membership Card"" for $35. Data mining + purchased loyalt"
Sumenn7063|HuffingtonPost|0.0|0.0|1.0|0.0|"RT @HuffingtonPost: Trevor Noah still can't figure out why Donald Trump calls China ""Jina"" https://t.co/qV216LQLMv https://t.co/lI5LkfdFpu"
Sumenn7063|m|0.0|0.0|1.0|0.0|"RT @HuffingtonPost: Trevor Noah still can't figure out why Donald Trump calls China ""Jina"" https://t.co/qV216LQLMv https://t.co/lI5LkfdFpu"
Gingersnap195|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
GlennLittle5|kausmickey|-0.6249|0.204|0.796|0.0|"RT @kausmickey: ""Trumps pick for Labor Secretary is perhaps the worst person imaginable for that role."" https://t.co/DiG5WsTVKU"
GlennLittle5|nationalreview|-0.6249|0.204|0.796|0.0|"RT @kausmickey: ""Trumps pick for Labor Secretary is perhaps the worst person imaginable for that role."" https://t.co/DiG5WsTVKU"
all10thingsNEWS|all10things|0.0|0.0|1.0|0.0|"Despite scientific consensus, Trump says nobody knows if climate change isrea https://t.co/pxlOljk0rJ"
kindnessNow16|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
LilushaLisa|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
MrAveryAvenue|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
medical_humor|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
medical_humor|thegatewaypundit|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
reanyc596|kylegriffin1|-0.5267|0.145|0.855|0.0|"RT @kylegriffin1: Watergate reporter Carl Bernstein: 'Nixon was nothing, in terms of lying, compared to what we've seen from Trump.' https:"
Sunshine2078|softwarnet|-0.8402|0.394|0.493|0.113|"@softwarnet @Eyes_of_justice the Dem outrage is real-Trump taxes ended up legal -DNC hacks exposed fraud, corruption, lies, &amp; spirit cooking"
Michelle82VHS|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
KevinARNG11BVet|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
asif_murdock|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
MPenny74|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
thiswaltz5|grumpyoldman418|0.5994|0.0|0.741|0.259|"RT @grumpyoldman418: Trump, Jr. Russians make up a pretty disproportionate cross-section of a lot of our assets,  https://t.co/ktNfyMSX9v"
thiswaltz5|linkis|0.5994|0.0|0.741|0.259|"RT @grumpyoldman418: Trump, Jr. Russians make up a pretty disproportionate cross-section of a lot of our assets,  https://t.co/ktNfyMSX9v"
BigBadBarb60|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
BigBadBarb60|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
nffc65|flyjawn|0.0|0.0|1.0|0.0|@flyjawn i would rather have snow than Trump
Rivera_Hugo|jnpaquet|0.34|0.0|0.897|0.103|RT @jnpaquet: Norwegian cartoonist Christian Bloom is creator of this cartoon of #Trump that has recently been shared on Twitter before cen
dogfriendlydude|Evan_McMullin|-0.1027|0.129|0.759|0.112|"RT @Evan_McMullin: Trump encouraged Russian subversion of our democracy then denied its occurrence despite CIA evidence, while preparing to"
hypnocoach183|MrJamesonNeat|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
hypnocoach183|t|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
ceili_woman|DLin71|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
ceili_woman|twitter|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
professorkck|twitter|-0.5267|0.134|0.866|0.0|This is who Trump and his team are. They crawled out of the right wing conspiracy sewer and will govern that way. D https://t.co/A647Dsgand
aboleyn|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
KyOgre_007|Jewrachi_007|0.0|0.0|1.0|0.0|"@Jewrachi_007 @GrouDonkey_007 One of these: Gary Johnson, Jill Stein, Donald Trump, Hillary Clinton"
benitah_summers|realjunsonchan|0.296|0.0|0.864|0.136|RT @realjunsonchan: Need to restore law and order in America #trump #maga #underdoges #americafirst https://t.co/m2R2CLxbo5
benitah_summers|twitter|0.296|0.0|0.864|0.136|RT @realjunsonchan: Need to restore law and order in America #trump #maga #underdoges #americafirst https://t.co/m2R2CLxbo5
DustinGiebel|JeffersonObama|0.0|0.0|1.0|0.0|RT @JeffersonObama: Trump never learned Russian until his 4th Bankruptcy #BoltonFalseFlagExcuses
MimiSteel|KeithOlbermann|0.0|0.0|1.0|0.0|RT @KeithOlbermann: CIA reveals how Russians ran a coup for Trump. From 10/14: the day Trump revealed he KNEW the Russians were doing it ht
NastierWoman|DavidYankovich|-0.1531|0.158|0.739|0.102|RT @DavidYankovich: My immediate goal is stopping Trump.Then we are going to end the GOP for their treason of the US by supporting enemie
klhgreen|BrentNYT|0.0|0.126|0.748|0.126|"RT @BrentNYT: The Russians hacked to support Trump - because they preferred a president they could manipulate, writes @nytopinion https://t"
klhgreen||0.0|0.126|0.748|0.126|"RT @BrentNYT: The Russians hacked to support Trump - because they preferred a president they could manipulate, writes @nytopinion https://t"
parker1313|jnpaquet|0.34|0.0|0.897|0.103|RT @jnpaquet: Norwegian cartoonist Christian Bloom is creator of this cartoon of #Trump that has recently been shared on Twitter before cen
jdprose|DLin71|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
jdprose|twitter|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
tata_colombia|twitter|0.0|0.0|1.0|0.0|"As te revuelques de la piedra, Trump (nada raro que l haga un tweet sobre esto) https://t.co/7BBdxAByx1"
other95|gollum1419_g|0.0|0.0|1.0|0.0|RT @gollum1419_g: Possible Trump Appointee Scrubs Facebook Post Fantasizing About Exterminating Muslims https://t.co/m3W7xL65AK #Resist #Tr
other95|rawstory|0.0|0.0|1.0|0.0|RT @gollum1419_g: Possible Trump Appointee Scrubs Facebook Post Fantasizing About Exterminating Muslims https://t.co/m3W7xL65AK #Resist #Tr
jyester55|activist360|0.0|0.0|1.0|0.0|RT @activist360: REPORT: Obsequious a**-kisser Trump's had his head up the colorectal cavities of Russian oligarchs for three decades https
lisbourne6|simon_schama|-0.5267|0.129|0.871|0.0|RT @simon_schama: Trump may just have been stupid enough to nominate for Sec of State the one person who turns the Russian election inquiry
_robertgraham|mattytalks|0.8479|0.0|0.638|0.362|"RT @mattytalks: In times like this it's important to speak truth to power. So I encourage everyone, write President Trump, tell him Beavis"
Momof4Lambs|ananavarro|-0.1027|0.136|0.746|0.118|"RT @ananavarro: Been off-line for hours vicariously suffering @MiamiDolphins' game...tell me, has Trump named Putin ""Special Advisor to the"
ric_m_martinez|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
DanceMyVoice|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
DanceMyVoice|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
DJTWATCHDOG|thetrumpwatchdog|0.0|0.0|1.0|0.0|Trump: US shouldnt be bound by one China Policy. https://t.co/IpO9basoSG
kvconstant|linkis|-0.4215|0.167|0.833|0.0|"Megyn Kelly says she fears reprisals for covering Trump, Breitbart News and the Alt-Right https://t.co/RpIE8dlRFd"
DebbiebB15|MelindaThinker|-0.4404|0.266|0.734|0.0|RT @MelindaThinker: Comey implicated in Trump Russia scandal https://t.co/OgZznjaH1f
DebbiebB15|bipartisanreport|-0.4404|0.266|0.734|0.0|RT @MelindaThinker: Comey implicated in Trump Russia scandal https://t.co/OgZznjaH1f
AliefofFaith|twitter|0.0|0.0|1.0|0.0|Obviously y'all from the part of Texas that voted for Trump https://t.co/sNe6CqWh4f
luckylucy061752|AndyOstroy|0.7003|0.126|0.504|0.37|RT @AndyOstroy: @ColMorrisDavis @JudgeJeanine @FoxNews Funny how these hypocrites prefer a draft-dodging coward over brave patriots like u
MLorance|politicususa|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
MLorance|twitter|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
soychilecl|soychile|0.0|0.0|1.0|0.0|"Donald Trump dijo que es ""ridcula"" la versin de que Rusia lo ayud a ganar https://t.co/63VDKILben https://t.co/ihN0QWojzS"
Jatapequara|chumbogrossomanaus|0.0|0.0|1.0|0.0|"Para Donald Trump reduzir as emisses de carbono prejudicam a competitividade global da Amrica e pergunta, ""Voc... https://t.co/GPQYqbyzHH"
Gojira007X|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
MDBeautyinOK|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Ohoura|BernieSanders|-0.3818|0.146|0.854|0.0|"RT @BernieSanders: Everyone who voted for Trump, who thought he'd defend working people, pay attention to the reality of what he's doing no"
PropersiDominic|LouDobbs|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
PropersiDominic|theconservativetreehouse|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
WTX11|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
smith_jeff999|MattOrtega|0.2732|0.0|0.851|0.149|"@MattOrtega Well, I don't know, just trying to be helpfulGlad for your trump site."
lindadoherty4|kurteichenwald|-0.5423|0.176|0.824|0.0|"RT @kurteichenwald: Fox/Cheney went nuts when found out Obama got intel briefings in writing, rather than read to him. But Trump no briefin"
TheSoundDefense|Anarky23|0.0|0.0|1.0|0.0|@Anarky23 Trump's ego is so fragile that a sneeze could shatter it
AllnattChris|realDonaldTrump|-0.7506|0.314|0.686|0.0|@realDonaldTrump @NBCNightlyNews @CNN Trump too weak to continue sanctions against Russia. In bed with the enemy.
cecemeddock|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
goldy_levy|raysr19|0.0|0.0|1.0|0.0|RT @raysr19: https://t.co/MnMVJMqO9J
goldy_levy|thegatewaypundit|0.0|0.0|1.0|0.0|RT @raysr19: https://t.co/MnMVJMqO9J
BuybyFelicia|jmaboshie|0.8573|0.165|0.482|0.354|"RT @jmaboshie: Im Vladimir, i stole the election for #Trump but I let Hillary win the popular vote. I forgot to rig that part. My bad. Won'"
rjennings333|dailymail|0.7579|0.0|0.698|0.302|Trump dismisses CIA claims that Russian hackers intervened to help him win election | Daily Mail Online https://t.co/3zat9Ru0zm
jonathankwonder|jnpaquet|0.34|0.0|0.897|0.103|RT @jnpaquet: Norwegian cartoonist Christian Bloom is creator of this cartoon of #Trump that has recently been shared on Twitter before cen
famdocparker1|SatPavanKaur|0.0|0.0|1.0|0.0|RT @SatPavanKaur: https://t.co/Cs1wDqRVcv Can the electoral college hold off on Trump until the country can figure what's going on. #TrumpL
famdocparker1|huffingtonpost|0.0|0.0|1.0|0.0|RT @SatPavanKaur: https://t.co/Cs1wDqRVcv Can the electoral college hold off on Trump until the country can figure what's going on. #TrumpL
RETTinol|instagram|0.0|0.0|1.0|0.0|foxnews's photo https://t.co/DwjXhBWIGy GO judge! TRUMP all the way!
TruthTeamOne|dem2119|0.4939|0.127|0.615|0.258|RT @dem2119: Dan Rather Just Called Out Fake Patriots Who Support Trumps Putin Romance In Viral Post - https://t.co/EIWDhA7hUu
TruthTeamOne|occupydemocrats|0.4939|0.127|0.615|0.258|RT @dem2119: Dan Rather Just Called Out Fake Patriots Who Support Trumps Putin Romance In Viral Post - https://t.co/EIWDhA7hUu
Beyoncelizer|beyonce|-0.6408|0.22|0.78|0.0|Race Baiter Beyonce Gets BAD News After Running Her Mouth at Trump - USA SUPREME... https://t.co/kjttjulZT0 https://t.co/vJ6EhvSFSM
cbl2|adamjohnsonNYC|-0.802|0.275|0.725|0.0|RT @adamjohnsonNYC: it was real news owning corporation Comcast--not fake news--that gave Trump a TV show after yrs of anti-black racism ht
unclesahm|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
unclesahm|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
deliamcmanus|mikeallen|0.2006|0.095|0.776|0.129|"RT @mikeallen: .@jimrutenberg column salutes @jaketapper: ""If only such moments could stop being so special and start being normal"" https:/"
deliamcmanus||0.2006|0.095|0.776|0.129|"RT @mikeallen: .@jimrutenberg column salutes @jaketapper: ""If only such moments could stop being so special and start being normal"" https:/"
BuffyMaxSFCA|tonyschwartz|0.7755|0.09|0.564|0.347|RT @tonyschwartz: Who cares that Trump doesn't believe Russians hacked Dems to elect him?Facts are indeed stubborn things &amp; the truth truly
lorac328|randyprine|-0.5859|0.147|0.853|0.0|RT @randyprine: NBC fires Billy Bush for listening to Trump brag about sexual assault yet Trump can Executive Produce a show on their netwo
ErickFernandez|charliek478|0.0|0.0|1.0|0.0|@charliek478 @PSheritaakkloh @Ckzoote https://t.co/O7Wrj6fdpW
ErickFernandez|politifact|0.0|0.0|1.0|0.0|@charliek478 @PSheritaakkloh @Ckzoote https://t.co/O7Wrj6fdpW
finscanes4life|CNNPolitics|0.4576|0.0|0.834|0.166|"RT @CNNPolitics: Israeli Prime Minister Benjamin Netanyahu: Donald Trump ""feels very warmly"" about Israel https://t.co/Vu0A4pgyce https://t"
finscanes4life|cnn|0.4576|0.0|0.834|0.166|"RT @CNNPolitics: Israeli Prime Minister Benjamin Netanyahu: Donald Trump ""feels very warmly"" about Israel https://t.co/Vu0A4pgyce https://t"
diegocosmelli|sciam|0.0|0.0|1.0|0.0|RT @sciam: An open letter from scientists to President-elect Trump on climate change https://t.co/A5DL4YVsuf https://t.co/WHKYXxg6Xb
diegocosmelli|blogs|0.0|0.0|1.0|0.0|RT @sciam: An open letter from scientists to President-elect Trump on climate change https://t.co/A5DL4YVsuf https://t.co/WHKYXxg6Xb
colbert_ed|twitter|0.0516|0.142|0.664|0.195|"A scary truth. New CIA will be filled with Trump loyalists &amp; disinformation specialists, nothing more than instrume https://t.co/fFYmqY6skb"
jmlilly|afreedma|0.1531|0.0|0.89|0.11|"RT @afreedma: Trump falsely claims that ""nobody knows"" if global warming is real https://t.co/RcgsNAPCPf"
jmlilly|mashable|0.1531|0.0|0.89|0.11|"RT @afreedma: Trump falsely claims that ""nobody knows"" if global warming is real https://t.co/RcgsNAPCPf"
huguetblanco|2016_Eleccion|0.0|0.0|1.0|0.0|"RT @2016_Eleccion: Biden: ""Trump hizo la campaa mas feroz que he visto"". https://t.co/QNFd06Dw1Q"
huguetblanco|twitter|0.0|0.0|1.0|0.0|"RT @2016_Eleccion: Biden: ""Trump hizo la campaa mas feroz que he visto"". https://t.co/QNFd06Dw1Q"
Paleoturkey|Trump_Supporter|-0.5423|0.412|0.588|0.0|@Trump_Supporter @c0nvey @YouTube It's a crime landslide.
ChrisSantana292|c0nvey|0.0|0.0|1.0|0.0|"""On Obamas watch, the economy generated 8.6 million net new jobs  or about... https://t.co/bI4hBdVpLD by #MarketWatch via @c0nvey"
ChrisSantana292|linkis|0.0|0.0|1.0|0.0|"""On Obamas watch, the economy generated 8.6 million net new jobs  or about... https://t.co/bI4hBdVpLD by #MarketWatch via @c0nvey"
kcarpe|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
chefdnel|StopPC101|0.0|0.0|1.0|0.0|@StopPC101 @realDonaldTrump Typical trump wuss can't handle the heat
ChavinhoMD|RT_com|-0.5256|0.152|0.848|0.0|RT @RT_com: #Hawking: Trumps victory &amp; Brexit come at the most dangerous time in the history of the human racehttps://t.co/wxW4JLIu2t
ymanesnah1|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
wendellshaw5|America_1st_|0.0|0.0|1.0|0.0|"RT @America_1st_: .@KellyannePolls: ""People who try to put Donald Trump in the conventional box are immediately and sorely disappointed."" h"
flyosity|tristanwalker|-0.5719|0.552|0.448|0.0|@tristanwalker Pathetic inconsistencies. https://t.co/ziogXd3mlx
flyosity|washingtonpost|-0.5719|0.552|0.448|0.0|@tristanwalker Pathetic inconsistencies. https://t.co/ziogXd3mlx
RR2969|Lrihendry|0.1275|0.113|0.756|0.13|RT @Lrihendry: While shopping 2day I overheard a conv with group saying isn't it great we can say Merry Christmas again &amp; not be afraid! WO
mrkisok|immigrant_legal|0.0|0.0|1.0|0.0|RT @immigrant_legal: Trump beat #NYTimes and #CNN at their own game https://t.co/0wdKh44NJe
mrkisok|twitter|0.0|0.0|1.0|0.0|RT @immigrant_legal: Trump beat #NYTimes and #CNN at their own game https://t.co/0wdKh44NJe
WishpathHealing|feministabulous|0.0|0.0|1.0|0.0|RT @feministabulous: i can't believe russia would hack the election after trump specifically asked them to https://t.co/V1dTFKOZOa
WishpathHealing|twitter|0.0|0.0|1.0|0.0|RT @feministabulous: i can't believe russia would hack the election after trump specifically asked them to https://t.co/V1dTFKOZOa
dukeblu85|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
dukeblu85|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
pharmalady|TearsInHeaven09|-0.5319|0.168|0.832|0.0|RT @TearsInHeaven09: LESSON:WHEN TRUMP TWEETS SOMETHING STUPIDHE IS TRYING TO MAKE YOU FORGETRUSSIA HACKED THE ELECTION FOR HIM
Seppie2727|sciam|0.0|0.0|1.0|0.0|RT @sciam: An open letter from scientists to President-elect Trump on climate change https://t.co/A5DL4YVsuf https://t.co/WHKYXxg6Xb
Seppie2727|blogs|0.0|0.0|1.0|0.0|RT @sciam: An open letter from scientists to President-elect Trump on climate change https://t.co/A5DL4YVsuf https://t.co/WHKYXxg6Xb
rew57|rtoberl|0.0|0.0|1.0|0.0|RT @rtoberl: John McCain doesn't know what to make of Trump's Russia hacking response https://t.co/2HyNt3zihL
rew57|linkis|0.0|0.0|1.0|0.0|RT @rtoberl: John McCain doesn't know what to make of Trump's Russia hacking response https://t.co/2HyNt3zihL
darrylwalter|businessinsider|-0.0772|0.098|0.902|0.0|Trump has shaken up decades of diplomacy with 4 phone calls #TrumpDanger  https://t.co/92FB0r31Cr https://t.co/T3d1jqVxPk
nancy73gg|LindaSuhler|0.0|0.0|1.0|0.0|RT @LindaSuhler: #PEOTUS Donald Trump &amp; Mike Pence #ThankYouTour2016 #PennsylvaniaHershey PAThurs 12/15 7 PM ET#MAGAReghttps://t.co
freemyheart31|childoflight4|-0.6597|0.302|0.554|0.144|"RT @childoflight4: 30% of Latinos (like me) LOVE Donald Trump yet these racist race baiting liars keep claiming its ""white people"" STOP THE"
AliasHere|dr_ashok_m|-0.5574|0.159|0.841|0.0|"RT @dr_ashok_m: It has to be #fakenews It cannot be Emails, foundation millions, #spiritcooking and Brazile cheating that caused @Hillary t"
DeLunaVintage|_dpaj|-0.296|0.239|0.638|0.122|"RT @_dpaj: Abortion Foes, Emboldened by Trump, Promise Onslaught of Tough Restrictions https://t.co/ZVzdFBvg7F ^NYTimes https://t.co/7dnh"
DeLunaVintage|nytimes|-0.296|0.239|0.638|0.122|"RT @_dpaj: Abortion Foes, Emboldened by Trump, Promise Onslaught of Tough Restrictions https://t.co/ZVzdFBvg7F ^NYTimes https://t.co/7dnh"
bebons101|CNNPolitics|0.0|0.0|1.0|0.0|"RT @CNNPolitics: Donald Trump: ""Nobody really knows"" if climate change is real https://t.co/BQ4z69MJJn https://t.co/Z9xI0BZ4Jt"
bebons101|cnn|0.0|0.0|1.0|0.0|"RT @CNNPolitics: Donald Trump: ""Nobody really knows"" if climate change is real https://t.co/BQ4z69MJJn https://t.co/Z9xI0BZ4Jt"
reanyc596|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
HubieDo|dailykos|0.0|0.0|1.0|0.0|Trump is laying the path for Democrats to reconsolidate the Blue Wall https://t.co/1jC5dp0o6o
jeffnews|dcexaminer|0.4019|0.0|0.778|0.222|"RT @dcexaminer: Allen West shares meme claiming Trump's defense secretary will ""exterminate"" Muslims https://t.co/oHZCB4uhtc https://t.co/D"
jeffnews|washingtonexaminer|0.4019|0.0|0.778|0.222|"RT @dcexaminer: Allen West shares meme claiming Trump's defense secretary will ""exterminate"" Muslims https://t.co/oHZCB4uhtc https://t.co/D"
marsam22reed|activist360|-0.5859|0.29|0.541|0.169|"RT @activist360: Trump admits his threat to lock up Clinton was just a prank to excite his hate-mongering, dirt dumb bigot base https://t.c"
marsam22reed||-0.5859|0.29|0.541|0.169|"RT @activist360: Trump admits his threat to lock up Clinton was just a prank to excite his hate-mongering, dirt dumb bigot base https://t.c"
Franield|kylegriffin1|-0.5267|0.145|0.855|0.0|"RT @kylegriffin1: Watergate reporter Carl Bernstein: 'Nixon was nothing, in terms of lying, compared to what we've seen from Trump.' https:"
LuciaBW15|P1e2h7Patrick|0.0516|0.0|0.93|0.07|RT @P1e2h7Patrick: Trump's cabinet serves purpose of legally tearing apart societal structure-Trump is authoritarian but foremost nihilist
FiveMeadows|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
jmingerson725|riotwomennn|0.296|0.0|0.879|0.121|"RT @riotwomennn: Russian Deputy Foreign Minister Sergei Ryabkov admits Russian gov ""maintained contacts"" w Trump during election  https://t"
jmingerson725||0.296|0.0|0.879|0.121|"RT @riotwomennn: Russian Deputy Foreign Minister Sergei Ryabkov admits Russian gov ""maintained contacts"" w Trump during election  https://t"
Tull007|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 7. Therefore, it could be a ""false flag"" operation by the Obama administration https://t.co/oRUPSkz7NV"
Tull007|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 7. Therefore, it could be a ""false flag"" operation by the Obama administration https://t.co/oRUPSkz7NV"
ProAssad|nytimesworld|0.0|0.0|1.0|0.0|"RT @nytimesworld: What if ""North Korea offers to Donald Trump that there is a lot of real estate that he can develop in North Korea""? https"
UT_MAZ|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
MikeSmithofABQ|rudepundit|-0.765|0.248|0.752|0.0|"RT @rudepundit: Maybe Trump is too dumb to understand that the word ""intelligence"" isn't meant as an insult to those being briefed."
Rajivkapoor2318|Newsmax|-0.6486|0.29|0.71|0.0|Michael Moore Plans to Protest at Trump Inauguration https://t.co/NLYMXzYmVq via @Newsmax Moore is an idiot
Rajivkapoor2318|newsmax|-0.6486|0.29|0.71|0.0|Michael Moore Plans to Protest at Trump Inauguration https://t.co/NLYMXzYmVq via @Newsmax Moore is an idiot
IngridWadsworth|Evan_McMullin|-0.5267|0.207|0.793|0.0|RT @Evan_McMullin: My Op-Ed in the NYTimes today: Trumps Threat to the Constitution https://t.co/6vNRZFaoxs
IngridWadsworth|nytimes|-0.5267|0.207|0.793|0.0|RT @Evan_McMullin: My Op-Ed in the NYTimes today: Trumps Threat to the Constitution https://t.co/6vNRZFaoxs
T_4an|realDonaldTrump|-0.8126|0.514|0.486|0.0|@realDonaldTrump @NBCNightlyNews @CNN pathetic Mr Trump you are pathetic.
Teleos|TeenVogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
Teleos|teenvogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
vickysue45|WeNeedTrump|0.0|0.0|1.0|0.0|RT @WeNeedTrump: Donald Trump and Mike Pence have the leadership we need to turn this country around. #MAGA https://t.co/pBokHtsx1y
vickysue45|twitter|0.0|0.0|1.0|0.0|RT @WeNeedTrump: Donald Trump and Mike Pence have the leadership we need to turn this country around. #MAGA https://t.co/pBokHtsx1y
OatesTuzzio|FoxNews|0.7925|0.0|0.713|0.287|@FoxNews @HillaryClinton she never said that. It's OK we know you've kissed up to Trump. U assume he's got 2 like one news outlet should b u
calnini|HamiltonElector|0.2298|0.123|0.757|0.12|"RT @HamiltonElector: Mr. Trump you are hardly a genius, no matter what Comrade Putin says.  We are smarter than you. We are #hamiltonelecto"
YaraM_A|JohnDelury|-0.7469|0.189|0.811|0.0|"RT @JohnDelury: Not to be alarmist, but when I asked what Beijing will do if Trump persists w Two China Policy, the answer was war https://"
YaraM_A||-0.7469|0.189|0.811|0.0|"RT @JohnDelury: Not to be alarmist, but when I asked what Beijing will do if Trump persists w Two China Policy, the answer was war https://"
EPICGOPFAIL|gerhadt_kreuz|-0.1027|0.142|0.733|0.125|"@gerhadt_kreuz @lisa5gk @skoobeedont Perhaps Russians/Trump cheated enough in Western PA + WI + MI 2 make this diff. turnout was good, tho"
miladysdewinter|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
tonic516|kurteichenwald|0.8607|0.0|0.677|0.323|"RT @kurteichenwald: GOP: Trump says doesnt need daily briefings cause he's so smart. So, u agree he is smarter than Reagan, who (like all o"
spaceyguys|helenmaryme|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
spaceyguys|twitter|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
Lermont|twitter|-0.5719|0.283|0.53|0.187|"Approaching a white Trump supporter &amp; assuming he's a racist, while assuming his black friend is not a racist is in https://t.co/Hgbz7nK5Vb"
BlueStateBob1|lillyslolly|-0.3724|0.131|0.869|0.0|"RT @lillyslolly: Donald Trump is 'not a loyal American', says former CIA operative and presidential candidate | The Independent https://t.c"
BlueStateBob1||-0.3724|0.131|0.869|0.0|"RT @lillyslolly: Donald Trump is 'not a loyal American', says former CIA operative and presidential candidate | The Independent https://t.c"
RachelK1967|funder|-0.2023|0.083|0.917|0.0|RT @funder: #TRUMPLEAKS:16 House Dems ask AG to investigate 25k bribe from Trump via Foundation for TrumpU#cnn #msnbc #AMJoy #cnnsotu #thi
WhosFibbing|_USAPolicalNewS|0.8971|0.0|0.479|0.521|RT @_USAPolicalNewS: Trumps BOLD NEW APPROACH to China is Brilliantly POWERFUL https://t.co/x23ieZoOX1 https://t.co/JzgNsgBkjZ
WhosFibbing|ilovemyfreedom|0.8971|0.0|0.479|0.521|RT @_USAPolicalNewS: Trumps BOLD NEW APPROACH to China is Brilliantly POWERFUL https://t.co/x23ieZoOX1 https://t.co/JzgNsgBkjZ
Tradekraft|foxnews|0.1511|0.0|0.923|0.077|"Kerry had ties to Iran, nothing was said !GOP senators challenge Trump on secretary of state prospect's Russia ties https://t.co/Uj7hIhzltO"
Joshua_A_Haney|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
Joshua_A_Haney|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
RobertSAdcock|2016Deplorables|0.5255|0.0|0.764|0.236|RT @2016Deplorables: Total respect! Army gives Trump his own jersey  #armynavy https://t.co/kYxR16XZX2
RobertSAdcock|twitter|0.5255|0.0|0.764|0.236|RT @2016Deplorables: Total respect! Army gives Trump his own jersey  #armynavy https://t.co/kYxR16XZX2
TheGrapesOfWisc|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
TheGrapesOfWisc|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
caitythekitty|kelseydarragh|-0.4404|0.176|0.758|0.066|RT @kelseydarragh: I keep acting like my problems r gunna b gone once 2016 is over but no Trump will b president and Im still gunna spend t
hanktastic1776|steph93065|0.0|0.0|1.0|0.0|RT @steph93065: To all the crazies following the Russian/Trump thing...Trump didn't give Russia enough uranium to nuke the entire world...
jaystebbins|Left_of_Texas|-0.4215|0.229|0.706|0.065|RT @Left_of_Texas: Dan Rather: Founding Fathers warned about a demagogue president backed by a foreign adversary - https://t.co/SIQRWZL8aV
jaystebbins|deadstate|-0.4215|0.229|0.706|0.065|RT @Left_of_Texas: Dan Rather: Founding Fathers warned about a demagogue president backed by a foreign adversary - https://t.co/SIQRWZL8aV
CharlieBrB|KeithOlbermann|0.0|0.0|1.0|0.0|RT @KeithOlbermann: CIA revealed Russia HAD tampered for Trump. From 10/14: when Trump revealed he knew they were doing it for him https://
CharlieBrB||0.0|0.0|1.0|0.0|RT @KeithOlbermann: CIA revealed Russia HAD tampered for Trump. From 10/14: when Trump revealed he knew they were doing it for him https://
TxMagnoliaLink|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
KarenCrow6|DailyCaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
KarenCrow6|dailycaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
dreamweaver1001|BrendanNyhan|0.0|0.0|1.0|0.0|RT @BrendanNyhan: Reminder: Trump has not disclosed finances that could reveal Russian ties &amp; could be enriched by them via businesses now
WendyJFluga28|BreitbartNews|0.2732|0.0|0.851|0.149|Report: Rick Perry on Trump's Energy Secretary Short List - Breitbart https://t.co/N7KInzo7wS via @BreitbartNews
WendyJFluga28|breitbart|0.2732|0.0|0.851|0.149|Report: Rick Perry on Trump's Energy Secretary Short List - Breitbart https://t.co/N7KInzo7wS via @BreitbartNews
brycedhowardfan|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
GonzaloWolfred|nytimes|0.0|0.0|1.0|0.0|Trump Suggests Using Bedrock China Policy as Bargaining Chip - New York Times https://t.co/5v1tEdRpdl
c_cathering|KeepAmerGr8|0.0|0.0|1.0|0.0|RT @KeepAmerGr8: Trump advisers with Russian ties https://t.co/n7szfoRLV6 via @msnbc
c_cathering|msnbc|0.0|0.0|1.0|0.0|RT @KeepAmerGr8: Trump advisers with Russian ties https://t.co/n7szfoRLV6 via @msnbc
vaveyla_t|nytimesworld|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
vaveyla_t|nytimes|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
ReclaimDawgs|vivelafra|-0.128|0.067|0.933|0.0|RT @vivelafra: Megyn Who? @TuckerCarlson is quickly becoming the biggest star on @FoxNews &amp; could dominate ratings for years to come. #Trum
JennyGardiner__|VoteHillary2016|0.0|0.0|1.0|0.0|"RT @VoteHillary2016: Trump's Secretary of State pick, @Exxon's @rex_tillerson, toasting Putin &amp; associates after signing lucrative deal. ht"
peanut96|nytimes|0.0|0.0|1.0|0.0|"""In Mr. Trump, the Russians had reason to see a malleable political novice..."" [can't wait to get T's tweet on this] https://t.co/NhpaB6qiKv"
JerseyStrong11|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
CountryLiberal|thedailybeast|0.0|0.0|1.0|0.0|"RT @thedailybeast: ""You voted for Donald Trump, thinking that he was on your side...Well, you got played."" - @JoyAnnReid: https://t.co/fKkb"
CountryLiberal|t|0.0|0.0|1.0|0.0|"RT @thedailybeast: ""You voted for Donald Trump, thinking that he was on your side...Well, you got played."" - @JoyAnnReid: https://t.co/fKkb"
tylerstone|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
tylerstone|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
gcamp4|twitter|0.0|0.0|1.0|0.0|This has been needed for so long and only Trump is the man for the job. The swamp draining will commence soon!! https://t.co/X1DbJ70Eb7
kh51048|LindaSuhler|-0.6239|0.23|0.678|0.092|@LindaSuhler Come 1/20/2017 cop killers will no longer have the support of the President. The real President will be after them. Go Trump!
NocturnalSu|THR|0.0|0.0|1.0|0.0|"RT @THR: ""Words have power. TV has power. My pen has power."" https://t.co/j7e4GjD3Pn"
NocturnalSu|hollywoodreporter|0.0|0.0|1.0|0.0|"RT @THR: ""Words have power. TV has power. My pen has power."" https://t.co/j7e4GjD3Pn"
dayadelreys|RuthHHopkins|0.5859|0.0|0.847|0.153|RT @RuthHHopkins: Russia helped Trump win. The CIA has confirmed this. The election is invalid. There's opinions &amp; there's facts. This is f
KandorKarteh|CaptainsLog2016|0.0|0.119|0.72|0.161|RT @CaptainsLog2016: Donald Trump said this word for wordOn national television&amp; now denies believing in any chance of Russia playing a
1775reaper|France4Hillary|-0.3612|0.128|0.872|0.0|"RT @France4Hillary: Given @CIA's evidence that Trump rigged the election with Russia, what should happen? #TrumPutingate #RussianHacking #L"
bani_amor|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
bani_amor||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
AlanAdrian3|V_of_Europe|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
AlanAdrian3|thegatewaypundit|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
LASmith3|NewtTrump|0.5267|0.0|0.861|0.139|"RT @NewtTrump: Newt explains Trump's MASTERFUL winning Twitter strategy ""If you don't give the media a rabbit to chase each day, they'll in"
havo1919|YouTube|-0.5423|0.289|0.597|0.114|The Truth About Fake News | Russia Hacked U.S. Election For Donald Trump? https://t.co/Y27qAuBbrM via @YouTube
havo1919|youtube|-0.5423|0.289|0.597|0.114|The Truth About Fake News | Russia Hacked U.S. Election For Donald Trump? https://t.co/Y27qAuBbrM via @YouTube
TheWestBay|Mtbkgrl|0.0|0.0|1.0|0.0|RT @Mtbkgrl: Trump licking Putin's ass...@realDonaldTrump#MAGA # FUCKINGPSYCOPATH https://t.co/0Ujl8f6HU4
TheWestBay|twitter|0.0|0.0|1.0|0.0|RT @Mtbkgrl: Trump licking Putin's ass...@realDonaldTrump#MAGA # FUCKINGPSYCOPATH https://t.co/0Ujl8f6HU4
LisaK4liberty|ed_hooley|-0.7213|0.209|0.791|0.0|"RT @ed_hooley: PUTIN DECLARES GEORGE SOROS IS A WANTED MAN DEAD OR ALIVEGeorge Soros's Home Address.136 Cantitoe St. Katonah, NY 10536#M"
OkcAllen|TheDemocrats|0.4939|0.0|0.802|0.198|RT @TheDemocrats: Trump has named: Anti-worker Labor SecretaryAnti-environment EPA admin.Anti-health care HHS SecretaryAnti-justice Att
mauree_b|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
mauree_b|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
SometimezY|noisey|-0.3612|0.143|0.857|0.0|Meet the Desi Artists Fighting Back Against Trump with Punk Rock and 'Post-Colonial Pop' - Noisey https://t.co/uR8cnn8KwP
Inked1BNA|SocialPowerOne1|0.3182|0.111|0.702|0.187|RT @SocialPowerOne1: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests https://t.co/Eghd6ic7s8
Inked1BNA|politicususa|0.3182|0.111|0.702|0.187|RT @SocialPowerOne1: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests https://t.co/Eghd6ic7s8
DaleMoss2|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: When Obama used Dijon mustard, Fox attackd him 4 not using yellow mustrd (true) Yet they shrug when Trump says doesnt n"
LFrady|FoxNews|0.5423|0.0|0.774|0.226|RT @FoxNews: Trump: We're Going to Start Saying 'Merry Christmas' Again https://t.co/rFmwtKQXIZ https://t.co/PexEqzNo9E
LFrady|insider|0.5423|0.0|0.774|0.226|RT @FoxNews: Trump: We're Going to Start Saying 'Merry Christmas' Again https://t.co/rFmwtKQXIZ https://t.co/PexEqzNo9E
hartsigns|jharlen00|-0.5719|0.198|0.802|0.0|"@jharlen00 @vandercyrus USA doesn't include the state trump lives in? your argument holds no water, she got 3 m more votes from AMERICANs"
centurionblog|GavinNewsom|-0.3089|0.101|0.899|0.0|RT @GavinNewsom: Trump's treating Russian interference in our election as partisan issue. This is not about political parties - our natl se
suesap1|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
ljanem|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
AhmadMunandar8|bt|0.0|0.0|1.0|0.0|Donald Trump varsler opgr med USA's et-Kina-politik - B.T. https://t.co/WlImlN65my
gjlos24|amjoyshow|0.0|0.0|1.0|0.0|RT @amjoyshow: Trump advisers with Russian ties https://t.co/hISlPTqQ2m via @amjoyshow
gjlos24|msnbc|0.0|0.0|1.0|0.0|RT @amjoyshow: Trump advisers with Russian ties https://t.co/hISlPTqQ2m via @amjoyshow
cocoabuttery|nbcnews|0.8316|0.109|0.461|0.431|Trump is too smart for daily briefings and too dumb to care about anything except himself  ha ha ha  https://t.co/V9j3ybHpFb
jocowboys87|JonRiley7|-0.0258|0.14|0.724|0.136|"RT @JonRiley7: ""Welcome to the Trump Administration, where climate change is fake and wrestling is real.""-- Trevor Noah"
bartbing71|medium|-0.7269|0.337|0.663|0.0|This is insane.  The US government is being taken over by conspiracy theorists.  https://t.co/kYwvWQkJ3O
Qrious123|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
Qrious123|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
DomAcconcia|AriMelber|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
DomAcconcia|t|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
jenbrunelle2|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
caroljdavy|JuddLegum|-0.3612|0.111|0.889|0.0|"RT @JuddLegum: 5. Bolton's evidence of this is that the CIA found evidence of Russian involvement, which he finds suspicious https://t.co/o"
caroljdavy|twitter|-0.3612|0.111|0.889|0.0|"RT @JuddLegum: 5. Bolton's evidence of this is that the CIA found evidence of Russian involvement, which he finds suspicious https://t.co/o"
princessmom122|eclecticbrotha|0.0|0.0|1.0|0.0|RT @eclecticbrotha: Three reasons Trump isn't taking intel briefings1. He can't read2. He wouldn't understand them if he could3. He pick
dwp1970|twitter|-0.7506|0.314|0.686|0.0|Student Threatened for Recording #triggered #Crybaby Teacher Who Called Trumps Election an Act of Terror - https://t.co/Vzc0SxZq8D
Presley48R|JewsChooseTrump|0.0516|0.11|0.714|0.176|"RT @JewsChooseTrump: #JewsChooseTrump Trump commits America to ""ensuring Israel maintains a qualitative military edge over all adversaries"""
smi26621356|CaptainKdog|-0.19|0.165|0.661|0.174|"RT @CaptainKdog: Trump first Pres. not only to BREAK campaign promises, but actively FIGHT AGAINST THEM. His Cabinet's history is OPPOSING"
cdo4Jesus|dayvarelat|0.128|0.0|0.914|0.086|RT @dayvarelat: Exclusive  First Day of Trumps Presidency: President-Elect Highlights Sacrifice of Americas Armed Forces at https://t
cdo4Jesus||0.128|0.0|0.914|0.086|RT @dayvarelat: Exclusive  First Day of Trumps Presidency: President-Elect Highlights Sacrifice of Americas Armed Forces at https://t
Who_R_U82|Mike_Padgett|0.0|0.0|1.0|0.0|RT @Mike_Padgett: '...most of what comes out of Trumps mouth is false...' https://t.co/cMGjY9tGS0
Who_R_U82|twitter|0.0|0.0|1.0|0.0|RT @Mike_Padgett: '...most of what comes out of Trumps mouth is false...' https://t.co/cMGjY9tGS0
jlmrbk|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
winged|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
jimstamant|andylassner|0.0431|0.123|0.713|0.163|RT @andylassner: Do NOT use this photo of Donald Trump. He does NOT like it. He told reporters he HATES it. Please RETWEET. https://t.c
jimstamant||0.0431|0.123|0.713|0.163|RT @andylassner: Do NOT use this photo of Donald Trump. He does NOT like it. He told reporters he HATES it. Please RETWEET. https://t.c
eileenpfeifer|RadioFreeTom|0.4767|0.0|0.876|0.124|"RT @RadioFreeTom: If HRC chose a SecState who ran an oil giant and got a medal from Putin, the GOPers defending Trump would re-convene the"
LisaToddSutton|SteveRattner|0.0|0.0|1.0|0.0|"RT @SteveRattner: With McCain and Graham opposed, will Tillerson (if he even gets nominated) be the first Trump pick to go down?"
SouthPawFaust|mikeoconnor123|-0.7906|0.32|0.68|0.0|"RT @mikeoconnor123: Press said  bi-partisan outrage if Trump challenged election, Then Hillary did just that.  Silence. Story on outrage is"
jjmplsmn|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
beemerjean|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
SonnyGirard|mikandynothem|0.3802|0.088|0.767|0.146|RT @mikandynothem: Ruth Bader Ginsburg said she would resign if Trump won. Hit the road lady! That will give Trump even more Conservatives
RoyClaflin|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
k_r_eckert|MicrotonalDan|0.0|0.0|1.0|0.0|RT @MicrotonalDan: FBI and CIA conclusions on Russia hacking don't line up https://t.co/vVrMgt5byV
k_r_eckert|cnn|0.0|0.0|1.0|0.0|RT @MicrotonalDan: FBI and CIA conclusions on Russia hacking don't line up https://t.co/vVrMgt5byV
sanesetti|HaikuVikingGal|-0.891|0.392|0.608|0.0|RT @HaikuVikingGal: Just a reminder that Donald Trump hates hates hates this photo of himself.  Do not retweet it. He hates it. https://t.c
sanesetti||-0.891|0.392|0.608|0.0|RT @HaikuVikingGal: Just a reminder that Donald Trump hates hates hates this photo of himself.  Do not retweet it. He hates it. https://t.c
danni_rie|JuddLegum|-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
danni_rie||-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
Sheljanz|ericgarland|-0.529|0.189|0.811|0.0|RT @ericgarland: The Russians didn't create Trump - only New York City and American gullibility could have done that.But they've got a SW
leeroyjenkins61|rickwells|0.6476|0.0|0.602|0.398|https://t.co/Gbg7OH5RwI  Energy Stocks will surely rise now! #MAGA #AmericaFirst #AltRight
GracefullyGray|yashar|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
GracefullyGray|twitter|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
Stphns|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
markevans08|MattAsherS|-0.1531|0.12|0.785|0.095|"RT @MattAsherS: @CheesbroV @markevans08 @MSNBC Sure, he has a right. Doesn't change fact that Trump criticism of intel &amp; media is irrespons"
irliteach|KenJennings|0.4404|0.0|0.884|0.116|RT @KenJennings: The Russians ABSOLUTELY have a sex tape of Trump and I just hope this ends without us having to watch any of it.
AnamikaMadad|HahnAmerica|-0.0572|0.06|0.94|0.0|RT @HahnAmerica: Why wouldn't Trump want a thorough bipartisan investigation of Russia hacking the DNC ? Why won't Trump release his taxes
efemmera|FeministaJones|-0.5106|0.18|0.82|0.0|RT @FeministaJones: Hey. I'm gonna be on c-span tomorrow morning talking about poverty in a Trump administration
ojhines2k|immigrant4trump|0.6588|0.0|0.82|0.18|RT @immigrant4trump: Video: Trump is going to Make America Great Again Regardless of the Color of your Skin! #Maga #Trump https://t.co/3aDj
ojhines2k|t|0.6588|0.0|0.82|0.18|RT @immigrant4trump: Video: Trump is going to Make America Great Again Regardless of the Color of your Skin! #Maga #Trump https://t.co/3aDj
dreamyswapnil|thehill|0.0|0.0|1.0|0.0|RT @thehill: Christie turned down several positions in Trump administration: reporthttps://t.co/Ff4dxZ0zkz https://t.co/LVefpPfmiC
dreamyswapnil|twitter|0.0|0.0|1.0|0.0|RT @thehill: Christie turned down several positions in Trump administration: reporthttps://t.co/Ff4dxZ0zkz https://t.co/LVefpPfmiC
wrahardian2|MAGAnNoHate|0.8555|0.0|0.567|0.433|@MAGAnNoHate @PioneerInvest Trump is the best for USA and the best for World
1975jetsfan4|BiasedGirl|0.0|0.0|1.0|0.0|RT @BiasedGirl: You know President-elect Trump is going to be tweeting about this... https://t.co/ZKymGISMXs
1975jetsfan4|twitter|0.0|0.0|1.0|0.0|RT @BiasedGirl: You know President-elect Trump is going to be tweeting about this... https://t.co/ZKymGISMXs
coolncalm3|MotherJones|-0.4215|0.135|0.865|0.0|@MotherJones @ToniJoseph14 not my sixties. If millenials keep protesting. It may mirror. But trump is in class by himself.
GingerAnnCazan|CaptainsLog2016|-0.5423|0.276|0.623|0.101|"RT @CaptainsLog2016: Dear @CanadaCan I book a 4 year stay in your country?I have no felonies, I pay taxes, and I didn't vote for Trump"
Napsterrific|NBCPolitics|0.0|0.0|1.0|0.0|RT @NBCPolitics: International students leery of Trump could cost U.S. billions https://t.co/AXrDnh6mFM
Napsterrific|nbcnews|0.0|0.0|1.0|0.0|RT @NBCPolitics: International students leery of Trump could cost U.S. billions https://t.co/AXrDnh6mFM
k3nnr|michelledozois|0.0|0.0|1.0|0.0|"RT @michelledozois: ""This is what Trump TV is."" https://t.co/p5777k3O80 https://t.co/CUeEKkysBd"
k3nnr|nytimes|0.0|0.0|1.0|0.0|"RT @michelledozois: ""This is what Trump TV is."" https://t.co/p5777k3O80 https://t.co/CUeEKkysBd"
adair_brion|yolandazavala7|0.0|0.0|1.0|0.0|RT @yolandazavala7: CIA Splinter Group Calls For Overthrow Of Trump Election https://t.co/qxAVFxYvA6 via @YouTube Watch for Constitutional
adair_brion|youtube|0.0|0.0|1.0|0.0|RT @yolandazavala7: CIA Splinter Group Calls For Overthrow Of Trump Election https://t.co/qxAVFxYvA6 via @YouTube Watch for Constitutional
ymanesnah1|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
SuburbanFemale|btiarao|0.0|0.0|1.0|0.0|"RT @btiarao: Wanna march for something? March for an end to voter suppression, which takes place in communities of color: https://t.co/N945"
SuburbanFemale|t|0.0|0.0|1.0|0.0|"RT @btiarao: Wanna march for something? March for an end to voter suppression, which takes place in communities of color: https://t.co/N945"
locvnguyen1|YouTube|-0.2263|0.203|0.638|0.159|OBAMA'S THREAT TO TURN THE MILITARY AGAINST TRUMP IS LIKE A CHIHUAHUA NI... https://t.co/4csIBAenwe via @YouTube
locvnguyen1|youtube|-0.2263|0.203|0.638|0.159|OBAMA'S THREAT TO TURN THE MILITARY AGAINST TRUMP IS LIKE A CHIHUAHUA NI... https://t.co/4csIBAenwe via @YouTube
tamiam71|MyPupVoted|-0.1391|0.223|0.577|0.2|@MyPupVoted @frankt370 Agree..haven't stopped Praying for God's hand to continue guiding Trump through..so sick of the corrupt left
CNCTBe|klookl|-0.3818|0.167|0.833|0.0|"Megyn Kelly Newt Gingrich FULL Interview Trump Polls , Fight Over Sexual Predator - https://t.co/DnYrszEMaN https://t.co/jqxsQgP0s4"
neonheretic|liamstack|0.0772|0.105|0.739|0.156|RT @liamstack: Now that Twitter has cracked down on the pro-Trump bots the top replies to @realDonaldTrump are mostly comedians mocking him
janet_yackle|WydenForOregon|0.0|0.0|1.0|0.0|I'm In: Let's Stand up to Trump! https://t.co/geK84EOOW4 via @WydenForOregon
janet_yackle|standtallforamerica|0.0|0.0|1.0|0.0|I'm In: Let's Stand up to Trump! https://t.co/geK84EOOW4 via @WydenForOregon
WBCBowie|twitter|-0.2235|0.112|0.888|0.0|This headline misrepresents what the article says.Your insinuating Trump is not hearing vital intelligence.This why https://t.co/ALCVyURxYM
bestpsychic4u|facebook|0.6483|0.117|0.566|0.317|Trump supporters: What was it that clinched your vote? The fake university? The less than charitable charity? The... https://t.co/PW3qfm4FiV
nanciemac|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
nanciemac|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
Cindy63306167|frankrichny|-0.1603|0.064|0.936|0.0|"RT @frankrichny: By holding back RNC emails, Putin didn't just help install Trump in White House but has means to blackmail GOP to do his b"
PIE20121|yashar|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
PIE20121|twitter|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
LSoudek|CaptainsLog2016|0.4767|0.0|0.807|0.193|RT @CaptainsLog2016: When someone tells you they believe Trump over the intelligence agencies https://t.co/uri6y47SkC
LSoudek|twitter|0.4767|0.0|0.807|0.193|RT @CaptainsLog2016: When someone tells you they believe Trump over the intelligence agencies https://t.co/uri6y47SkC
TidyStucco_com|bloomberg|-0.34|0.194|0.806|0.0|Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/9oxwgbjV3k https://t.co/3qRtPfPaJw
rdanielkelemen|TheEconomist|0.34|0.119|0.693|0.188|"RT @TheEconomist: Republicans are denying that Russias authoritarian, anti-American government wanted Mr Trump to win https://t.co/WGgzEMk"
rdanielkelemen|t|0.34|0.119|0.693|0.188|"RT @TheEconomist: Republicans are denying that Russias authoritarian, anti-American government wanted Mr Trump to win https://t.co/WGgzEMk"
jyester55|abctweet100|-0.4404|0.206|0.7|0.093|RT @abctweet100: Trump Ignores National Security Facts When It Doesn't Suit Him #USA We Are Screwed #HamiltonElectors YOUR OBLIGATION IS TO
dredeyedick|youtube|-0.1779|0.116|0.884|0.0|Six More Women Come Forward Accusing Presumptive PEOTUS Donald Trump of #SexualAssault https://t.co/QbOTOREqey #ElectoralCollege
rachmanworks|CNBC|0.0|0.0|1.0|0.0|"RT @CNBC: Trump says U.S. not necessarily bound by ""one China"" policy https://t.co/hkRFMZLkxO"
rachmanworks|cnbc|0.0|0.0|1.0|0.0|"RT @CNBC: Trump says U.S. not necessarily bound by ""one China"" policy https://t.co/hkRFMZLkxO"
gitanalatina07|ananavarro|-0.1027|0.136|0.746|0.118|"RT @ananavarro: Been off-line for hours vicariously suffering @MiamiDolphins' game...tell me, has Trump named Putin ""Special Advisor to the"
axgueca|UniPolitica|0.0|0.0|1.0|0.0|"RT @UniPolitica: Trump vuelve a desdear la informacin de la CIA sobre el posible hackeo de Rusia: ""Es ridculo"" https://t.co/VZdWNu5xKr h"
axgueca|univision|0.0|0.0|1.0|0.0|"RT @UniPolitica: Trump vuelve a desdear la informacin de la CIA sobre el posible hackeo de Rusia: ""Es ridculo"" https://t.co/VZdWNu5xKr h"
RosalesRosina|ezlusztig|0.0|0.0|1.0|0.0|"RT @ezlusztig: I've noticed on the far right that this term ""false flag"" is getting thrown at anything that seems to compromise Trump."
tlvrp_russia|rt|0.0|0.0|1.0|0.0|#Moscow #SaintPetersburg Netanyahu has about 5 ideas for Trump to undo Iran nuclear deal https://t.co/HNYb7x9hpC
linda_wed1|funder|-0.6808|0.286|0.714|0.0|RT @funder: Criminal Complaint being filed on Donald Trump-for TREASON-for involvement w/Russia hack #news#TrumpLeaks #russiahacking #wat
roqchrisy|Trump_Commander|-0.7003|0.279|0.721|0.0|RT @Trump_Commander: VIDEO : Trump Responds to Crazy Liberals Russian Conspiracy Theories Every Week Its Something New https://t.co/LUZr
roqchrisy|t|-0.7003|0.279|0.721|0.0|RT @Trump_Commander: VIDEO : Trump Responds to Crazy Liberals Russian Conspiracy Theories Every Week Its Something New https://t.co/LUZr
PortugalLiving|BrendanNyhan|-0.7579|0.28|0.669|0.05|"@BrendanNyhan If Trump swears to defend constitution ""against enemies foreign ..."" would this lie constitute a High Crime and Misdemeanor?"
claytonorama|rabihalameddine|0.0|0.0|1.0|0.0|RT @rabihalameddine: I'm way too old to try and understand people who voted for Trump. https://t.co/SQU1hyfS6e
claytonorama|twitter|0.0|0.0|1.0|0.0|RT @rabihalameddine: I'm way too old to try and understand people who voted for Trump. https://t.co/SQU1hyfS6e
LisaQuake|twitter|-0.5255|0.236|0.764|0.0|"Broken machines, Russian hackers, voter suppression...how can anyone call #Trump President?! https://t.co/cao8QPaYaf"
Gav_Kumar|tech|0.7845|0.0|0.653|0.347|US intelligence analysts conclude that Russia helped Trump win the 2016 elections https://t.co/tuAIdxQcUF https://t.co/pvCLNXJm07 Tech
LozierJeannine|StuPolitics|0.6113|0.052|0.709|0.239|RT @StuPolitics: Why on earth are the Trump folks so defensive about this?  He won the election. Their defensiveness is laughable and ridic
jennifer4nm|kurteichenwald|0.5574|0.0|0.847|0.153|"RT @kurteichenwald: If Trump started getting praise 4  appointments from ISIS, do you think Fox News would start running stories about how"
Teresa_H_|LouDobbs|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
Teresa_H_|theconservativetreehouse|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
DoreeeV|TeamTrump|0.0|0.0|1.0|0.0|RT @TeamTrump: How the market looks one month after a Trump win:'biggest 1-month S&amp;P 500 rally in its 93 yrs of existence'https://t
Mainiac1820New|twitter|0.0772|0.131|0.679|0.19|"WSJ https://t.co/xnnVG1D9DZ his recent attacks on corporate America, Trump said: I want us to make good deals fo https://t.co/mF7f5u85uK"
davecfields|AntTheIcon|0.4515|0.141|0.617|0.242|RT @AntTheIcon: worst 2 teams? 49ers with a BLM QB and the BROWNS. best record? the AMERICAN conference PATRIOTS whose QB publicly supports
Tespis|c0nvey|0.0|0.0|1.0|0.0|'#Tolerant' city #making #Trump kids' lives horrible... https://t.co/w7cwBkdq2K by #StCyrlyMe2 via @c0nvey
Tespis|linkis|0.0|0.0|1.0|0.0|'#Tolerant' city #making #Trump kids' lives horrible... https://t.co/w7cwBkdq2K by #StCyrlyMe2 via @c0nvey
MHPspeechballon|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
badaboom100|RonaldKlain|0.0|0.0|1.0|0.0|"RT @RonaldKlain: This is not ""normal:""  Today, Trump tweeted cancellation of a contract, employing thousands, after reading that Boeing had"
i_vamshi|forbes|0.0|0.0|1.0|0.0|Donald Trump's $100 Million Private Jet Features Gold-Plated (Nearly) Everything https://t.co/XNHjA3LagE https://t.co/mG991AXXdw
Brock4Liberty|jnpaquet|0.34|0.0|0.897|0.103|RT @jnpaquet: Norwegian cartoonist Christian Bloom is creator of this cartoon of #Trump that has recently been shared on Twitter before cen
SitnokGlobal|markets|-0.128|0.209|0.613|0.178|RT @markets: Mexico's creditworthiness is under threat because of Trump https://t.co/pBXDVRoUpX https://t.co/mihf7BVDbp
SitnokGlobal|bloomberg|-0.128|0.209|0.613|0.178|RT @markets: Mexico's creditworthiness is under threat because of Trump https://t.co/pBXDVRoUpX https://t.co/mihf7BVDbp
JeannieM0625|ValkyrieHanna7|0.3724|0.0|0.825|0.175|@ValkyrieHanna7 U didnt listen 2 her bcuz ur #MSM didnt report it Shame on u.https://t.co/VnMIUBBr5L
rcivmares88|sarahkendzior|0.0|0.0|1.0|0.0|RT @sarahkendzior: Here is what Harry Reid wrote to James Comey about Trump-Russia collusion. US citizens deserve to know. https://t.co/lsI
rcivmares88|t|0.0|0.0|1.0|0.0|RT @sarahkendzior: Here is what Harry Reid wrote to James Comey about Trump-Russia collusion. US citizens deserve to know. https://t.co/lsI
Andrianamik|ed_hooley|-0.7213|0.209|0.791|0.0|"RT @ed_hooley: PUTIN DECLARES GEORGE SOROS IS A WANTED MAN DEAD OR ALIVEGeorge Soros's Home Address.136 Cantitoe St. Katonah, NY 10536#M"
Tommywa|le_Parisien|0.0|0.0|1.0|0.0|RT @le_Parisien: Etats-Unis : Trump : Je ne veux pas que la Chine me dicte ce que je dois faire https://t.co/GI2gGn9boc
Tommywa|l|0.0|0.0|1.0|0.0|RT @le_Parisien: Etats-Unis : Trump : Je ne veux pas que la Chine me dicte ce que je dois faire https://t.co/GI2gGn9boc
DCCorners|nytimes|0.1779|0.173|0.602|0.226|Can Congress End Donald Trump's Conflict of Interest Exemption? https://t.co/A24X9Kg7gX
ujhsteacher|randyprine|0.3612|0.079|0.753|0.168|"RT @randyprine: Instead of vilifying the CIA, Trump should release his taxes to prove that Russia has no incentive for helping him be elect"
TamarGranor|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
thejoecool|asterios|-0.2023|0.114|0.886|0.0|RT @asterios: [11 women accuse Trump of assault]They're shills.[CIA says Russia interfered]No way.[Podesta mentions pizza]THEY'RE
daxis_gaming|RamonaCallender|-0.2023|0.122|0.878|0.0|@RamonaCallender strange then why did trump say some parts will be fenced not wall
THETRUT80439582|truth-ng|0.5319|0.0|0.762|0.238|"COME OVER TO NIGERIA AND HELP US, FAYOSE URGES TRUMP. https://t.co/W61ydKrgqH https://t.co/uuFHtOZA75"
dervishmandala|historyinflicks|-0.3612|0.106|0.894|0.0|RT @historyinflicks: Trump in Nov: the election could be rigged. i might not concede.Dems in Dec: change dot org petition asking the Deep
DebbiebB15|DailyNewsBin|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
DebbiebB15|palmerreport|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
wklei1|randyprine|0.3612|0.079|0.753|0.168|"RT @randyprine: Instead of vilifying the CIA, Trump should release his taxes to prove that Russia has no incentive for helping him be elect"
JoinerMari|funder|-0.4404|0.17|0.83|0.0|RT @funder: #TrumpLeaks: Pam Bondi-Florida AG who took bribe to drop #trumpu cases-mtg w/Trump today for admin post #payforplay #msnbc #cnn
Koryatstirling|Esquire|-0.25|0.118|0.882|0.0|Trump's 'America-First' Plan Is Already Going Up in Flames https://t.co/p5dMEASwVy via @Esquire @realDonaldTrump screws his voters
Koryatstirling|esquire|-0.25|0.118|0.882|0.0|Trump's 'America-First' Plan Is Already Going Up in Flames https://t.co/p5dMEASwVy via @Esquire @realDonaldTrump screws his voters
nellss20|TeenVogue|0.4019|0.115|0.691|0.194|"RT @TeenVogue: .@realDonaldTrump is gaslighting America and undermining the very foundation of our freedom, by @laurenduca https://t.co/lxH"
nellss20|t|0.4019|0.115|0.691|0.194|"RT @TeenVogue: .@realDonaldTrump is gaslighting America and undermining the very foundation of our freedom, by @laurenduca https://t.co/lxH"
HonkyTonkNights|hannity|0.0|0.0|1.0|0.0|"Despite Boeing's Claims, Trump's $4 Billion Price Tag For New Air Force Ones Is Accurate https://t.co/oUVJdlGiwL"
PresidentBoyd|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
PresidentBoyd||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
RayeAlbright|VOANews|0.5859|0.0|0.769|0.231|RT @VOANews: Possible Tillerson Choice for US Top Diplomat Raises Questions of Corporate vs National Interest https://t.co/D2S6uKjyTH https
RayeAlbright|voanews|0.5859|0.0|0.769|0.231|RT @VOANews: Possible Tillerson Choice for US Top Diplomat Raises Questions of Corporate vs National Interest https://t.co/D2S6uKjyTH https
koons_rob|SenJohnMcCain|0.5499|0.0|0.843|0.157|@SenJohnMcCain @FaceTheNation @CBSNews Russia did zero to sway this election.   The media swayed it but interestingly they swayed to Trump
NSaneMotivation|thehill|0.0|0.0|1.0|0.0|"RT @thehill: Trump consulting lawyers on adding Ivanka, Jared Kushner to administrationhttps://t.co/xta6rFJUoh https://t.co/wfZ3aSrxbK"
NSaneMotivation|twitter|0.0|0.0|1.0|0.0|"RT @thehill: Trump consulting lawyers on adding Ivanka, Jared Kushner to administrationhttps://t.co/xta6rFJUoh https://t.co/wfZ3aSrxbK"
azenkova2|wikileaks|-0.4021|0.153|0.763|0.084|"@wikileaks I'm GOD'S Voice! God says:""I'll change all your Elite on Earth! TRUMP is only the BEGINNING! LIBERALS will DISAPPEAR soon!God"""
moskaezul|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
adammizelle|saladinahmed|-0.3818|0.11|0.89|0.0|RT @saladinahmed: there are ten thousand reasons that anyone with any shred of decency should fight trump.'he doesn't listen to the CIA'
AndreMinn|expansion|0.0|0.0|1.0|0.0|Walmart desestima a Trump al anunciar inversiones en Mxico? https://t.co/YNvDToQWm8 https://t.co/nxZUwsMuFk
TalLouis111|Will_Bunch|-0.7149|0.239|0.761|0.0|"RT @Will_Bunch: Worse than Watergate? Russia hacking is massive cloud over Trump presidency, and America. What caused this big mess? https:"
EmotioNerd|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
iAm_KJayy|QveenTee6|0.0772|0.0|0.925|0.075|RT @QveenTee6: trump should make it mandatory for everyone to take lessons on HOW TO TEXT BACK
brettbeletz|ashleyn1cole|-0.296|0.109|0.891|0.0|RT @ashleyn1cole: Everyone Trump has picked wants to dismantle the agency they will be running. That's it. No punchline.
Archin2014|Joyce_Karam|-0.8176|0.309|0.691|0.0|RT @Joyce_Karam: There's an attack on Church in Egypt;Terror in Istanbul; ISIS took Palmyra; CIA alarm on Russia.But #Trump is attacking NB
ChatterTNN|WhitevsBIackTwt|-0.0191|0.097|0.903|0.0|RT @WhitevsBIackTwt: hillary and trump will never reach this level https://t.co/goPD3NSnmC
ChatterTNN|vine|-0.0191|0.097|0.903|0.0|RT @WhitevsBIackTwt: hillary and trump will never reach this level https://t.co/goPD3NSnmC
Uberskiper|RepAdamSchiff|0.1027|0.12|0.741|0.139|RT @RepAdamSchiff: Conflicts of interest Trump will bring into oval office are unprecedented. #ActLikeAPresident &amp; divest completely. @nyti
Bayathread|margaretcho|0.5859|0.0|0.703|0.297|@margaretcho follow @RachelleHodgs for brilliant graphing of Trump word salads.
NetCatNews|twitter|0.2023|0.0|0.833|0.167|#news #summary: top tech leaders to meet with  #trump https://t.co/lIlnK4UzeT
PeterBacon5|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
roqchrisy|asamjulian|0.8934|0.0|0.592|0.408|"RT @asamjulian: Not that the popular vote matters, but Trump won the popular vote by 2+ million in 49 states. https://t.co/OMS2M0flDu"
roqchrisy|twitter|0.8934|0.0|0.592|0.408|"RT @asamjulian: Not that the popular vote matters, but Trump won the popular vote by 2+ million in 49 states. https://t.co/OMS2M0flDu"
MrJamesJoint|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/TEGHqhLpZN https://t.co"
MrJamesJoint|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/TEGHqhLpZN https://t.co"
micah_gideon|slate|-0.5267|0.167|0.833|0.0|"Had anyone reading this heard of the ""Pizza Sex Conspiracy"" before learning its promoters are on Trump's team?https://t.co/yQplIGGDb6"
DeathsHead725|DJTrump45|0.0|0.0|1.0|0.0|RT @DJTrump45: The #Trump45 Daily! https://t.co/im4eFFJLE7 #trump
DeathsHead725|paper|0.0|0.0|1.0|0.0|RT @DJTrump45: The #Trump45 Daily! https://t.co/im4eFFJLE7 #trump
vishesh81|FT|-0.7964|0.323|0.677|0.0|RT @FT: The dangers of Donald Trumps coming boom. @edwardGLuce on the temptation to undermine Fed and scapegoat China https://t.co/BeRziwB
vishesh81|t|-0.7964|0.323|0.677|0.0|RT @FT: The dangers of Donald Trumps coming boom. @edwardGLuce on the temptation to undermine Fed and scapegoat China https://t.co/BeRziwB
raemadema|Suntimes|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
raemadema|chicago|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
Positividad3|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: The Big Oil Allies and Beltway Insiders Leading Trumps Department of the Interior  and How to by @JamesCTobias https://
Positividad3||0.0|0.0|1.0|0.0|RT @starfirst: The Big Oil Allies and Beltway Insiders Leading Trumps Department of the Interior  and How to by @JamesCTobias https://
AlbertWarner|ScottAdamsSays|0.7249|0.0|0.568|0.432|@ScottAdamsSays Trump blogs as AUDIOBOOK with you reading please. thanks!!!
Unicorn688|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
Unicorn688|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
rowemichael|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
realtimb|jnpaquet|0.34|0.0|0.897|0.103|RT @jnpaquet: Norwegian cartoonist Christian Bloom is creator of this cartoon of #Trump that has recently been shared on Twitter before cen
E__R__O|frankrichny|-0.1603|0.064|0.936|0.0|"RT @frankrichny: By holding back RNC emails, Putin didn't just help install Trump in White House but has means to blackmail GOP to do his b"
tabishch|forbes|0.0|0.0|1.0|0.0|Donald Trump's $100 Million Private Jet Features Gold-Plated (Nearly) Everything https://t.co/6B7zB9MMH1 via #Tashify.com #MavoTV.com
aurojm|SinEmbargoMX|-0.5423|0.163|0.837|0.0|"RT @SinEmbargoMX: Heisenberg, de Breaking Bad, candidato a dirigir la DEA con Donald Trump. Al menos en SNL https://t.co/Ie6GsIWj2X https:/"
aurojm|sinembargo|-0.5423|0.163|0.837|0.0|"RT @SinEmbargoMX: Heisenberg, de Breaking Bad, candidato a dirigir la DEA con Donald Trump. Al menos en SNL https://t.co/Ie6GsIWj2X https:/"
Djs12377|TheDemocrats|0.5514|0.0|0.818|0.182|RT @TheDemocrats: Are you:- A woman?- Under 26?Do you:- Have a pre-existing condition?- Live?- Breathe?Obamacare helps you. Don't le
klknott|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
Eric_111|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
KenBerry611|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
KenBerry611|change|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
huggafop|Slate|0.0|0.0|1.0|0.0|RT @Slate: Exxon Mobil's CEO is frontrunner to be Trump's Secretary of State. Here's what the company's been up to on his watch https://t.c
huggafop||0.0|0.0|1.0|0.0|RT @Slate: Exxon Mobil's CEO is frontrunner to be Trump's Secretary of State. Here's what the company's been up to on his watch https://t.c
matygarcia|PolticsNewz|0.0|0.0|1.0|0.0|RT @PolticsNewz: Russia's head of foreign affairs applaud's Trump's secretary of State pick https://t.co/YChWVoCG9f https://t.co/1jcqOir1FI
matygarcia|route|0.0|0.0|1.0|0.0|RT @PolticsNewz: Russia's head of foreign affairs applaud's Trump's secretary of State pick https://t.co/YChWVoCG9f https://t.co/1jcqOir1FI
bigbill_ontw|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
Amertunesucre|davebernstein|-0.296|0.131|0.784|0.086|RT @davebernstein:  CALL TO ACTION: Please call the DOJ at # below &amp; tell them you are outraged re: Russian interference to elect Donald T
RT_CNN|money|-0.6249|0.24|0.76|0.0|#news #trump #hillary #election #syria These are the world's worst tax havens https://t.co/aw7brunObW https://t.co/izKdgtFgKL
ajitsinghpundir|buyindian|-0.6597|0.226|0.726|0.048|"RT @buyindian: If anything 'laughable and ridiculous' is poor American people who believe in US Democracy, When Trump selling US.  https://"
ajitsinghpundir||-0.6597|0.226|0.726|0.048|"RT @buyindian: If anything 'laughable and ridiculous' is poor American people who believe in US Democracy, When Trump selling US.  https://"
KimBL13|vivelafra|-0.6486|0.194|0.806|0.0|"RT @vivelafra: BIG 6: After criminally colluding with his opponent for 18 months, MSM is now trying to suggest #Trump had an unfair advanta"
FoolishlyHigh|BernieSanders|-0.3818|0.146|0.854|0.0|"RT @BernieSanders: Everyone who voted for Trump, who thought he'd defend working people, pay attention to the reality of what he's doing no"
tonic516|funder|-0.2023|0.083|0.917|0.0|RT @funder: #TRUMPLEAKS:16 House Dems ask AG to investigate 25k bribe from Trump via Foundation for TrumpU#cnn #msnbc #AMJoy #cnnsotu #thi
shirl47char|ed_hooley|-0.7213|0.209|0.791|0.0|"RT @ed_hooley: PUTIN DECLARES GEORGE SOROS IS A WANTED MAN DEAD OR ALIVEGeorge Soros's Home Address.136 Cantitoe St. Katonah, NY 10536#M"
Lindalizer|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Lindalizer||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
ManceKathy|thehill|0.0|0.0|1.0|0.0|https://t.co/PYE9Yh62dM
anneh1313|SenSanders|0.4767|0.08|0.691|0.229|"RT @SenSanders: I challenge Mr. Trump to tell the American people he'll keep his promises and veto cuts to Social Security, Medicare and Me"
instinctnaturel|RepAdamSchiff|0.1027|0.12|0.741|0.139|RT @RepAdamSchiff: Conflicts of interest Trump will bring into oval office are unprecedented. #ActLikeAPresident &amp; divest completely. @nyti
Tull007|JuddLegum|0.5979|0.0|0.811|0.189|"RT @JuddLegum: 6. According to Bolton, Russians are so good at hacking they would never leave evidence that US intel could detect https://t"
Tull007||0.5979|0.0|0.811|0.189|"RT @JuddLegum: 6. According to Bolton, Russians are so good at hacking they would never leave evidence that US intel could detect https://t"
tanyachambers81|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
KTowns17|RawStory|0.0|0.0|1.0|0.0|RT @RawStory: Possible Trump appointee scrubs Facebook post after fantasizing about exterminating Muslims https://t.co/bW4F2tc0OL https:/
KTowns17|rawstory|0.0|0.0|1.0|0.0|RT @RawStory: Possible Trump appointee scrubs Facebook post after fantasizing about exterminating Muslims https://t.co/bW4F2tc0OL https:/
TLee5T|simonhelberg|0.8126|0.0|0.657|0.343|RT @simonhelberg: cool just go on instinct I'm sure there's not much to this whole president thing oh my god help https://t.co/uqnX4BatOq
TLee5T|medium|0.8126|0.0|0.657|0.343|RT @simonhelberg: cool just go on instinct I'm sure there's not much to this whole president thing oh my god help https://t.co/uqnX4BatOq
Left_of_Labor|Broelman|0.0|0.0|1.0|0.0|RT @Broelman: Trumpushka #trump #trumpadministration #Trumpageddon #auspol https://t.co/Y7ovMvujKl
Left_of_Labor|twitter|0.0|0.0|1.0|0.0|RT @Broelman: Trumpushka #trump #trumpadministration #Trumpageddon #auspol https://t.co/Y7ovMvujKl
SinsBeggar|realDonaldTrump's|0.4588|0.0|0.727|0.273|A #limerick fer @realDonaldTrump's favorite picture.#NotMyPresident #PresidentBitchBoy #Trump #TrumpLeaks https://t.co/5lk45lkUUA
SinsBeggar|twitter|0.4588|0.0|0.727|0.273|A #limerick fer @realDonaldTrump's favorite picture.#NotMyPresident #PresidentBitchBoy #Trump #TrumpLeaks https://t.co/5lk45lkUUA
carolinesreflex|c0nvey|0.0|0.0|1.0|0.0|It took me seconds to realise that it's trump's face. https://t.co/rdlnmBupgk by #Scorpio_A7 via @c0nvey
carolinesreflex|linkis|0.0|0.0|1.0|0.0|It took me seconds to realise that it's trump's face. https://t.co/rdlnmBupgk by #Scorpio_A7 via @c0nvey
worldnews_net|theglobeandmail|-0.0516|0.066|0.934|0.0|"Rex Tillerson, Trumps likely secretary of state, is a life-long oil man who backs Keystone https://t.co/no62MB7qpL #Globe #Mail #news"
aramiscat|funder|0.0|0.0|1.0|0.0|RT @funder: Donald Trump called me David &amp; himself Goliath.I don't think he knows how that ended#TrumpIsBeingInvestigated!#TrumpLeaks
WhoIsDEF|KenJennings|0.4404|0.0|0.884|0.116|RT @KenJennings: The Russians ABSOLUTELY have a sex tape of Trump and I just hope this ends without us having to watch any of it.
caroljdavy|JuddLegum|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
caroljdavy|t|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
cbendik79|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
cbendik79||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
THRGlobal|realDonaldTrump|0.1027|0.206|0.619|0.175|Wanda Chairman and China's Richest Man Warns @realDonaldTrump About Blocking Chinese Investment in U.S. https://t.co/r2ILXC4MQI
THRGlobal|twitter|0.1027|0.206|0.619|0.175|Wanda Chairman and China's Richest Man Warns @realDonaldTrump About Blocking Chinese Investment in U.S. https://t.co/r2ILXC4MQI
JimRousch|realDonaldTrump|-0.4767|0.22|0.78|0.0|To state the obvious: @realDonaldTrump is wrong.  https://t.co/RB97k3xIuS by #puppymnkey via @c0nvey
JimRousch|linkis|-0.4767|0.22|0.78|0.0|To state the obvious: @realDonaldTrump is wrong.  https://t.co/RB97k3xIuS by #puppymnkey via @c0nvey
murph7041|0ryuge|-0.1838|0.138|0.752|0.11|@0ryuge @RobotShlomo @jahimes @cliffschecter too bad a minority of ppl cannot see how stupid trump is and the con job being done.
kmkinnaird|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
AtomicShock2012|jacobmathews|-0.2732|0.211|0.655|0.135|RT @jacobmathews: @SenJohnMcCain cyber attacks been happening for years. Why the urgency now?  Is  that because your foe Trump won Presiden
Perpetual_Now|gant1014|-0.2808|0.164|0.723|0.113|"RT @gant1014: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/pJ2y2vUpSR via @Bipartisan Re"
Perpetual_Now|bipartisanreport|-0.2808|0.164|0.723|0.113|"RT @gant1014: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/pJ2y2vUpSR via @Bipartisan Re"
JulioGautreaux|FoxNews|0.5848|0.0|0.774|0.226|"RT @FoxNews: President-elect @realDonaldTrump: ""We're going to start saying 'Merry Christmas' again!"" https://t.co/rFmwtKzmkp https://t.co/"
JulioGautreaux|insider|0.5848|0.0|0.774|0.226|"RT @FoxNews: President-elect @realDonaldTrump: ""We're going to start saying 'Merry Christmas' again!"" https://t.co/rFmwtKzmkp https://t.co/"
ChuckOlson5|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
ChuckOlson5||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
DeborahRacona|MikePenceVP|0.091|0.097|0.791|0.112|"RT @MikePenceVP: No, Donald Trump isn't going to attack gay rights, women's rights, religious minoritys. Because he isn't practicing radi"
Shanny_resqchi|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
Shanny_resqchi|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
_Carolina_Man_|MarkDice|0.8146|0.065|0.65|0.285|@MarkDice #MSM self-destructed in 2016 to our delight! What we suspected became oh so apparent! Much fun seeing Trump smack the #FakeNews!
tlvrp_russia|therussophile|0.25|0.0|0.882|0.118|"#Moscow #SaintPetersburg Trumps personality unprecedented, vision of new world order yet to be seen  Kissinger https://t.co/0yIgG8gHOM"
Iraclestic|Giants|0.2263|0.185|0.573|0.242|Wow even Donald Trump Hates Erick Flowers performance #NYGvsDAL @Giants https://t.co/GBY4ertjtk
Iraclestic|twitter|0.2263|0.185|0.573|0.242|Wow even Donald Trump Hates Erick Flowers performance #NYGvsDAL @Giants https://t.co/GBY4ertjtk
BitcoinBuddhist|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
BitcoinBuddhist|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
RNRoxx|JeffreyGuterman|0.5267|0.085|0.698|0.217|"RT @JeffreyGuterman: . @LizWahl: ""The goal of Russian media is to undermine faith in our institutions and now they've succeeded in hacking"
audispeak|DeanLeh|-0.5413|0.163|0.837|0.0|RT @DeanLeh: Draining the swamp? TRUMP IS the swamp &amp; has surrounded himself with very scary swamp creatures. #ThanksYouIgnorantTrumpVoters
Fails_us|forbes|0.0|0.0|1.0|0.0|Donald Trump's $100 Million Private Jet Features Gold-Plated (Nearly) Everything https://t.co/Oz75HmIYfK https://t.co/qDn8XkfoiM
NewsInTweetsCom|newsintweets|0.0|0.0|1.0|0.0|Huffington Post: Most Americans dont think Trump should have to sell his companies to be president https://t.co/vinSnHtrb5 #NewsInTweets
KilianJulianus|washingtontimes|0.0|0.169|0.663|0.169|"Donald Trump-Tsai Ing-wen phone call raises hopes, fears in Taiwan - Washington Times https://t.co/4Y1dwZAgQW"
tedreally|yashar|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
tedreally|twitter|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
grandpooba5440|riotwomennn|-0.3724|0.113|0.887|0.0|RT @riotwomennn: Former CIA operative &amp; House GOP aide Evan McMullin: 'Trump is not a loyal American'  Are you listening Electors?  https:/
grandpooba5440||-0.3724|0.113|0.887|0.0|RT @riotwomennn: Former CIA operative &amp; House GOP aide Evan McMullin: 'Trump is not a loyal American'  Are you listening Electors?  https:/
MarkGisler|greenhousenyt|-0.2732|0.095|0.905|0.0|RT @greenhousenyt: Unions underestimated Trump's appeal to the working classNow he &amp; GOP lawmakers will seek to hobble laborMy Story: htt
loregraf|ActualidadRT|0.0|0.0|1.0|0.0|RT @ActualidadRT: Trump critica a la CIA por acusar a Rusia https://t.co/LvSjecKd7e
loregraf|actualidad|0.0|0.0|1.0|0.0|RT @ActualidadRT: Trump critica a la CIA por acusar a Rusia https://t.co/LvSjecKd7e
HWOZONE|alexjonesshows|-0.4019|0.162|0.838|0.0|RT @alexjonesshows: Trump dismisses the CIAs claim it has evidence Russians hacked the election https://t.co/BlIQajTzOd
HWOZONE|alexjonespodcast|-0.4019|0.162|0.838|0.0|RT @alexjonesshows: Trump dismisses the CIAs claim it has evidence Russians hacked the election https://t.co/BlIQajTzOd
SusanaCanabal|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
Andy_J_Crawford|KeithOlbermann|0.0|0.0|1.0|0.0|RT @KeithOlbermann: CIA revealed Russia HAD tampered for Trump. From 10/14: that time Trump revealed he knew they were doing it for him htt
THECROWSTWEET|Bikers4Trump|-0.4588|0.149|0.785|0.066|@Bikers4Trump @Quoimio @CeciliaFrances4 @Bikers_4_Trump Hear ya bro. If intentions are solid don't sweat the small shit &amp; just do your thing
DonetaKP|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
jlseaback|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
hollyoptix|NewYorker|0.2263|0.109|0.727|0.164|RT @NewYorker: .@BorowitzReport: Poll: Americans Favor Keeping Air Force One and Cancelling Trump https://t.co/MGQdWsegjM
hollyoptix|newyorker|0.2263|0.109|0.727|0.164|RT @NewYorker: .@BorowitzReport: Poll: Americans Favor Keeping Air Force One and Cancelling Trump https://t.co/MGQdWsegjM
ChrisRosche|FrankLuntz|0.0|0.0|1.0|0.0|"RT @FrankLuntz: ""How do you brief a president who refuses to believe what you tell him?""https://t.co/W2vLESP6l2"
ChrisRosche|politico|0.0|0.0|1.0|0.0|"RT @FrankLuntz: ""How do you brief a president who refuses to believe what you tell him?""https://t.co/W2vLESP6l2"
TallDarkNotUgly|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
MagnusDahlgren|TIME|0.0|0.0|1.0|0.0|RT @TIME: Meet the voters who helped put Donald Trump in the White House #TIMEPOY https://t.co/i4fJn9EQqA
MagnusDahlgren|time|0.0|0.0|1.0|0.0|RT @TIME: Meet the voters who helped put Donald Trump in the White House #TIMEPOY https://t.co/i4fJn9EQqA
NetCatNews|twitter|0.0|0.0|1.0|0.0|"#news #summary:  #trump says  #wall  #street journal doesn't ""understand  #business"" https://t.co/MMvFsfZYnw"
djsandwiches|Suntimes|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
djsandwiches|chicago|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
bdascholten|wsj|0.34|0.088|0.772|0.14|Always someone to blame. Worked to win; will it work to govern and lead? Trump Fuels Rift With CIA Over Russian Hack https://t.co/PV3jtEcLs4
tlvrp_russia|therussophile|0.0|0.0|1.0|0.0|#Moscow #SaintPetersburg PHOTOS: Rogue One Premiere Targeted by Pro-Trump Street Artist https://t.co/GLCDX4FH5h
janewicjane|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
janewicjane|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
mypostdemise|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
GlennF|liamstack|0.0772|0.105|0.739|0.156|RT @liamstack: Now that Twitter has cracked down on the pro-Trump bots the top replies to @realDonaldTrump are mostly comedians mocking him
JeffersonObama|JPMendelson|0.6908|0.0|0.759|0.241|RT @JPMendelson: Trump eats bacon cheeseburgers and other fast food regularly. At 70. Giving him to 90 is generous. https://t.co/vOdsCArBDB
JeffersonObama|twitter|0.6908|0.0|0.759|0.241|RT @JPMendelson: Trump eats bacon cheeseburgers and other fast food regularly. At 70. Giving him to 90 is generous. https://t.co/vOdsCArBDB
busdog|BernieSanders|-0.1531|0.122|0.778|0.1|RT @BernieSanders: Donald Trump is a pathological liar.  We need the help of the American people to build a movement of millions who are fo
tlvrp_russia|therussophile|0.6369|0.0|0.634|0.366|#Moscow #SaintPetersburg Watch: Trump Greeted With Cheers at Army-Navy Game https://t.co/emlLJhqlFC
WallaceGreene|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
WallaceGreene||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
teakinrj|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
teakinrj||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
robtmackinnon|JuddLegum|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
robtmackinnon|t|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
uchiyama4949|jp|0.0|0.0|1.0|0.0| |  https://t.co/RmeIIHJR3s _(*c
Deteacherintell|npr|0.0|0.0|1.0|0.0|FACT CHECK: Trump Claims A 'Massive Landslide Victory'  But History Differs https://t.co/L0FsMLFJD0
jocowboys87|laureldavilacpa|0.0|0.0|1.0|0.0|RT @laureldavilacpa: #ImStillNotOver Before the election the Senate was briefed by the CIA of #RussianHackers electioneering for Trump - an
RayMaso75618253|JonRiley7|-0.0258|0.14|0.724|0.136|"RT @JonRiley7: ""Welcome to the Trump Administration, where climate change is fake and wrestling is real.""-- Trevor Noah"
TheJoshLoweShow|independent|0.2607|0.127|0.695|0.179|Donald Trump says he doesn't need daily intelligence briefings as President because he's 'smart' - fantastic https://t.co/OHK1Be2H51
baloo035|Evan_McMullin|-0.1027|0.129|0.759|0.112|"RT @Evan_McMullin: Trump encouraged Russian subversion of our democracy then denied its occurrence despite CIA evidence, while preparing to"
tlvrp_russia|therussophile|0.0|0.0|1.0|0.0|"#Moscow #SaintPetersburg Reid Wont Go Away: Russian Involvement In Election A Hanging Chad 1,000 Times Over, Tr https://t.co/3txTIn42Ms"
cphillip3|NBCPolitics|0.0|0.0|1.0|0.0|RT @NBCPolitics: International students leery of Trump could cost U.S. billions https://t.co/AXrDnh6mFM
cphillip3|nbcnews|0.0|0.0|1.0|0.0|RT @NBCPolitics: International students leery of Trump could cost U.S. billions https://t.co/AXrDnh6mFM
LisaMoraitis1|dem2119|0.4939|0.127|0.615|0.258|RT @dem2119: Dan Rather Just Called Out Fake Patriots Who Support Trumps Putin Romance In Viral Post - https://t.co/EIWDhA7hUu
LisaMoraitis1|occupydemocrats|0.4939|0.127|0.615|0.258|RT @dem2119: Dan Rather Just Called Out Fake Patriots Who Support Trumps Putin Romance In Viral Post - https://t.co/EIWDhA7hUu
paraluman_uk|DrEstella|0.0|0.0|1.0|0.0|"RT @DrEstella: Senator #HarryRead asks CIA to lie to @realDonaldTrump ""Give Trump ""Fake"" INTEL BRIEFINGS!""  #SundayMorning #WeareTrump #Tru"
washumom|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
cheapskare|starfirst|-0.6908|0.213|0.787|0.0|RT @starfirst: Donald Trump and the Republican's leaders are guilty of treason. They're  traitors  of the very soil they stand on they are
BershodM|occupydemocrats|-0.4939|0.211|0.789|0.0|SNL Just Destroyed Trumps Narcissism With This Hillarious Through Donalds Eyes Skit - https://t.co/TFgKtSLCoN
keithahodges|merica_man84|0.3612|0.0|0.815|0.185|"@merica_man84 @CNN Bannon White Nazi=Russian ,Sessions Putin wants a trump dictatorship like Russia"
OLSXWatching|medium|-0.765|0.423|0.577|0.0|Trumps lies have a purpose. They are an assault on democracy https://t.co/9TZWk5TNve
brixtondoyle|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
brixtondoyle|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
DucinniAnthony|YouTube|-0.5904|0.204|0.796|0.0|INSIDER: TRUMP TO PULL PLUG ON FAKE CLIMATE CHANGE AGENDA MAKE US ENERGY... https://t.co/d3FX6193RH via @YouTube
DucinniAnthony|youtube|-0.5904|0.204|0.796|0.0|INSIDER: TRUMP TO PULL PLUG ON FAKE CLIMATE CHANGE AGENDA MAKE US ENERGY... https://t.co/d3FX6193RH via @YouTube
LMoelhauser|KeithOlbermann|0.5362|0.0|0.886|0.114|RT @KeithOlbermann: We now know what the Russians did for Trump. Next: what is he doing for them? From 9/28: Is he loyal to the US? 9/28 ht
linda_wed1|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: Trump: 'Nobody really knows' if #ClimateChange is real. Um... Apart from every scientist who works on the subject?! Idi
amicuss|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
rbean14620|WillBlackWriter|0.3182|0.0|0.897|0.103|RT @WillBlackWriter: Please tweet and ask your followers to tweet this Vine of Donald Trump asking Russia to hack Clinton. #Treasonhttps
goldy_levy|JackPosobiec|-0.2168|0.161|0.719|0.12|RT @JackPosobiec: You mean like how you worked to defeat Trump's nomination? How'd that go again? https://t.co/3petpHwFvj
goldy_levy|twitter|-0.2168|0.161|0.719|0.12|RT @JackPosobiec: You mean like how you worked to defeat Trump's nomination? How'd that go again? https://t.co/3petpHwFvj
tlvrp_russia|therussophile|-0.2263|0.137|0.863|0.0|"#Moscow #SaintPetersburg California Elector Files Lawsuit, Joins Movement to Find Trump Alternative https://t.co/TiFYjSa0jv"
rohit0761|forbes|0.0|0.0|1.0|0.0|Donald Trump's $100 Million Private Jet Features Gold-Plated (Nearly) Everything https://t.co/4SzGMZJab0 https://t.co/yWi3PMO4gn
pgarcialujan|nymag|0.3567|0.159|0.607|0.234|I've never loved this beautiful blue bubble quite as much as I do now. https://t.co/YURioSLvvu
esteban_nieves|YourAnonCentral|-0.4939|0.144|0.856|0.0|"RT @YourAnonCentral: Steal this: Open Call for mobilization against the inauguration of Donald #Trump on January 20, 2017 #DisruptJ20  http"
Dystopianna|ezlusztig|0.0|0.0|1.0|0.0|RT @ezlusztig: Source: https://t.co/dh3On46A0t
Dystopianna|theguardian|0.0|0.0|1.0|0.0|RT @ezlusztig: Source: https://t.co/dh3On46A0t
alanpdx|JoyAnnReid|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
alanpdx|twitter|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
StandingsNYC|MarkRuffalo|0.4767|0.0|0.823|0.177|"RT @MarkRuffalo: Why does Putin want Trump Pres? $500 billion opportunity for Exxon, Russia in Trump cabinet pick | MSNBC #ExxonKnew  https"
marineshamus|NewssTrump|0.5267|0.0|0.825|0.175|"RT @NewssTrump: VIDEO : Democrat Congresswoman Praises Trump, Says Obama Admin is Funding Al-Qaeda and ISIS https://t.co/HiekEB3VEx https:/"
marineshamus|truthfeed|0.5267|0.0|0.825|0.175|"RT @NewssTrump: VIDEO : Democrat Congresswoman Praises Trump, Says Obama Admin is Funding Al-Qaeda and ISIS https://t.co/HiekEB3VEx https:/"
rdnktk|MrDane1982|0.0|0.0|1.0|0.0|"RT @MrDane1982: Part of the CIA investigation should be a deeper look into Donald Trump finances while releasing his tax returns, his deep"
IceMarinos|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
Pixelfish|ScottMadin|-0.4939|0.165|0.752|0.083|"RT @ScottMadin: I'm so old I remember when ""Donald Trump"" was a clich joke about how fucked up New York was in the '80s"
SandraPitts14|funder|-0.2023|0.083|0.917|0.0|RT @funder: #TRUMPLEAKS:16 House Dems ask AG to investigate 25k bribe from Trump via Foundation for TrumpU#cnn #msnbc #AMJoy #cnnsotu #thi
pinklady404|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
Rickeyleetw|ed_hooley|-0.7213|0.209|0.791|0.0|"RT @ed_hooley: PUTIN DECLARES GEORGE SOROS IS A WANTED MAN DEAD OR ALIVEGeorge Soros's Home Address.136 Cantitoe St. Katonah, NY 10536#M"
srauer20|leahmcelrath|0.5719|0.0|0.812|0.188|@leahmcelrath @blogdiva @brownblaze if he turns on trump I WILL take pleasure in it...so little of that nowadays
richminer|rstevens|0.3818|0.105|0.673|0.222|"RT @rstevens: Hate to admit it, but I support Trumps choice of Cigarette Smoking Man for Surgeon General https://t.co/QDvLTsca85"
richminer|twitter|0.3818|0.105|0.673|0.222|"RT @rstevens: Hate to admit it, but I support Trumps choice of Cigarette Smoking Man for Surgeon General https://t.co/QDvLTsca85"
LaurelSnyder|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
MrsESK|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
SC_Ropp|Khanoisseur|-0.4404|0.139|0.861|0.0|"RT @Khanoisseur: While US media snoozed, Financial Times did reported on how dirty money flowed into Trump @SamSanderson123 @summerbrennan"
DeathsHead725|mitchellvii|0.7914|0.108|0.56|0.332|"RT @mitchellvii: I would not be surprised if Russia favored Trump winning.  After 8 years, they didn't want another idiot running America."
OuelletteVicky|France4Hillary|-0.4514|0.217|0.616|0.167|RT @France4Hillary: It makes me SO SICK to see that Trump is lying about the Russian help he received to win the election. MAN UP &amp; TELL TH
danknapp76|MichaelGaree|-0.5267|0.204|0.739|0.057|"RT @MichaelGaree: Something comrade Trump's inner circle might want to consider: If he's charged with treason, guess who becomes co-conspir"
sewingsandra|America_1st_|0.8248|0.0|0.708|0.292|"RT @America_1st_: CW: ""The thing that impressed me was that Trump is always comfortable in own skin, but now he was comfortable being the P"
JimmyMak1|trumpwallnow|0.8689|0.073|0.541|0.385|@trumpwallnow Ha yes we've already discussed that. Trump won. America lost. Including you. But you probably trust Russia over US too right?
maddie142519|cmwarnerstl|0.4019|0.0|0.856|0.144|RT @cmwarnerstl: @Playfulimp @VABVOX @BernieSanders Yes he was.  The Devine - Manafort connection is the Bernie - Trump connection.
Tull007|JuddLegum|-0.3612|0.111|0.889|0.0|"RT @JuddLegum: 5. Bolton's evidence of this is that the CIA found evidence of Russian involvement, which he finds suspicious https://t.co/o"
Tull007|twitter|-0.3612|0.111|0.889|0.0|"RT @JuddLegum: 5. Bolton's evidence of this is that the CIA found evidence of Russian involvement, which he finds suspicious https://t.co/o"
JBucknoff|washingtonpost|-0.3612|0.152|0.848|0.0|#Trump shows his ignorance by falsely claiming nobody really knows if #climatechange is real. https://t.co/7t6WKxLNJZ
MarlaJ101|JonHutson|-0.3724|0.203|0.797|0.0|RT @JonHutson: Repeat: Donald Trump is not a loyal American. #resist https://t.co/s9j6SE1Mif
MarlaJ101|twitter|-0.3724|0.203|0.797|0.0|RT @JonHutson: Repeat: Donald Trump is not a loyal American. #resist https://t.co/s9j6SE1Mif
Dainesi1616|HirokoTabuchi|0.4215|0.0|0.859|0.141|RT @HirokoTabuchi: Not true. The $50 billion will come from a previously announced $100 billion investment fund. https://t.co/vLpqF9x72K @r
Dainesi1616|cnbc|0.4215|0.0|0.859|0.141|RT @HirokoTabuchi: Not true. The $50 billion will come from a previously announced $100 billion investment fund. https://t.co/vLpqF9x72K @r
394Hunter|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
ABCBTom|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
ABCBTom|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
0463diamond|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
Zhape|rdlaing|-0.8271|0.34|0.584|0.076|"RT @rdlaing: My take:Clinton: Let me explain about the emails   Press: Liar liar liar   Trump: I lie, its what I do.   Press: Ok"
su_z_t|"DavidYankovich)So,"|0.2732|0.0|0.861|0.139|"Retweeted David Yankovich (@DavidYankovich):So, Donald Trump has committed treason... This is a moment for... https://t.co/poGGUFz1Ds"
su_z_t|facebook|0.2732|0.0|0.861|0.139|"Retweeted David Yankovich (@DavidYankovich):So, Donald Trump has committed treason... This is a moment for... https://t.co/poGGUFz1Ds"
Latersbaby_28|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
LKuehn4|kurteichenwald|0.4215|0.0|0.877|0.123|RT @kurteichenwald: .@SenJohnMcCain - briefed on intel - say on air that he knows evidence of Russian interference and its true. Trump team
nickmjimenez|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
tip1665|mikandynothem|0.4404|0.0|0.868|0.132|RT @mikandynothem: President-elect Trump hasn't even taken Office yet and he's already showing himself to be a better President than Obama.
paintbygretzky|IMPL0RABLE|0.0|0.0|1.0|0.0|RT @IMPL0RABLE: #TheResistance Hamilton electorsThis makes 10California elector joins anti-Trump #ElectoralCollege push https://t.co/aV
paintbygretzky|t|0.0|0.0|1.0|0.0|RT @IMPL0RABLE: #TheResistance Hamilton electorsThis makes 10California elector joins anti-Trump #ElectoralCollege push https://t.co/aV
Kashinka|MtnMD|-0.2023|0.087|0.913|0.0|"RT @MtnMD: RT @PhiKapMom: Ryan, McConnell, Comey-&gt;any GOP involved in covering up Russian involvement in election for Trump needs charged i"
ChristianRep|BIZPACReview|0.8221|0.0|0.691|0.309|"RT @BIZPACReview: Total respect! Troops show their love for Trump at Army-Navy game; check out the video, photos https://t.co/Mv7RDPbKLg"
ChristianRep|bizpacreview|0.8221|0.0|0.691|0.309|"RT @BIZPACReview: Total respect! Troops show their love for Trump at Army-Navy game; check out the video, photos https://t.co/Mv7RDPbKLg"
stanhopekevin|starfirst|0.1779|0.076|0.812|0.112|"RT @starfirst: John McCain, Lindsey Graham join with Democrats to demand answers on Russias pro-Trump hacking https://t.co/4RUAylYaQG via"
stanhopekevin|dailynewsbin|0.1779|0.076|0.812|0.112|"RT @starfirst: John McCain, Lindsey Graham join with Democrats to demand answers on Russias pro-Trump hacking https://t.co/4RUAylYaQG via"
slidewinding|funder|0.8176|0.0|0.706|0.294|"RT @funder: Breaking: Ku Klux Klan parades in Roxboro, NC celebrating Trump win #cnn #msnbc #ncpol #amjoy #antitrump #trumpleaks https://t."
slidewinding||0.8176|0.0|0.706|0.294|"RT @funder: Breaking: Ku Klux Klan parades in Roxboro, NC celebrating Trump win #cnn #msnbc #ncpol #amjoy #antitrump #trumpleaks https://t."
amandablount2|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
amandablount2|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
AngryJackRabbit|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
StephenRBeck1|CNN|-0.8088|0.216|0.784|0.0|@CNN @CNNOpinion SO STUPID CNN!!  Putin would much rather walk all over hillary any day than try to push Trump around.  THINK ABOUT THAT!!!!
ReeeVamped718|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: When Obama used Dijon mustard, Fox attackd him 4 not using yellow mustrd (true) Yet they shrug when Trump says doesnt n"
jadedsquirrel|helenmaryme|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
jadedsquirrel|twitter|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
anibal__lopez|TooLitConcerts|-0.4404|0.209|0.791|0.0|RT @TooLitConcerts: Schoolboy Q on stage about how much he hates Trump  https://t.co/Ko6Q6W92gD
anibal__lopez|twitter|-0.4404|0.209|0.791|0.0|RT @TooLitConcerts: Schoolboy Q on stage about how much he hates Trump  https://t.co/Ko6Q6W92gD
transgarrus|meganamram|0.0|0.0|1.0|0.0|RT @meganamram: Real question: does Trump believe in object permanence
HoosierMum|thenation|0.0258|0.15|0.694|0.156|"RT @thenation: Democrats Should Fight All of Trumps Nominees. Yes, All of Them. https://t.co/gJZxnQv7fQ"
HoosierMum|thenation|0.0258|0.15|0.694|0.156|"RT @thenation: Democrats Should Fight All of Trumps Nominees. Yes, All of Them. https://t.co/gJZxnQv7fQ"
jitzkow52|nytopinion|0.0|0.0|1.0|0.0|RT @nytopinion: Why would President-elect Trump object to a thorough bipartisan probe into Russian meddling? https://t.co/zDopY4Hcs0 https:
jitzkow52|nytimes|0.0|0.0|1.0|0.0|RT @nytopinion: Why would President-elect Trump object to a thorough bipartisan probe into Russian meddling? https://t.co/zDopY4Hcs0 https:
j_b_trey|twitter|0.4404|0.104|0.677|0.219|I disagree. 60 million donkeys voted for Trump and all the GOP henchmen. I hope this will motivate voters for next https://t.co/UgGwUQqS1c
queenreee|SkepticPugilist|0.0|0.0|1.0|0.0|RT @SkepticPugilist: Just to put this into context: Trump wants to jail people who burn the American flag for longer than Brock Turner got
RohanElessar|realDonaldTrump|0.6597|0.0|0.779|0.221|"Trump says ""he's smart"" so he doesn't need briefings everyday. @realDonaldTrump If you have to tell people you're smart, you're not."
Chambord22|AWill83192048|-0.8126|0.345|0.576|0.079|RT @AWill83192048: @MrDane1982 Bernie: Its all riggedTrump: Its all rigged biglyAmericans: Hell yeah it was rigged for Trump.BS &amp; DT: c
bbdevices|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
bbdevices||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
CarmenRaye|JoyAnnReid|0.4019|0.0|0.828|0.172|RT @JoyAnnReid: They are the party of Trump. All previous monikers are extinct. https://t.co/f92tTxy7z8
CarmenRaye|twitter|0.4019|0.0|0.828|0.172|RT @JoyAnnReid: They are the party of Trump. All previous monikers are extinct. https://t.co/f92tTxy7z8
Markus03121966|SimonWDC|-0.5849|0.159|0.841|0.0|RT @SimonWDC: The most troubling aspect of the Russia story is how much Trump has embraced Putin's worldview.  More here: https://t.co/kqUE
Markus03121966|t|-0.5849|0.159|0.841|0.0|RT @SimonWDC: The most troubling aspect of the Russia story is how much Trump has embraced Putin's worldview.  More here: https://t.co/kqUE
giddeygirl|nobby15|0.0|0.0|1.0|0.0|"RT @nobby15: Republicans to launch wide-ranging probe of Russia election hacking, despite Trump's stance https://t.co/3HjcQc2Ucb via @Radio"
giddeygirl|abc|0.0|0.0|1.0|0.0|"RT @nobby15: Republicans to launch wide-ranging probe of Russia election hacking, despite Trump's stance https://t.co/3HjcQc2Ucb via @Radio"
mimix3|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
mnoxides|FoxNews|-0.1779|0.124|0.876|0.0|RT @FoxNews: .@JudgeJeanine Slams Obama: 'Why Are You Obsessed With Russia?' https://t.co/96TVMVqFc9 https://t.co/WkwW8sYfbg
mnoxides|insider|-0.1779|0.124|0.876|0.0|RT @FoxNews: .@JudgeJeanine Slams Obama: 'Why Are You Obsessed With Russia?' https://t.co/96TVMVqFc9 https://t.co/WkwW8sYfbg
bulldogfinance|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
SamLo91|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
ujhsteacher|randyprine|0.0|0.0|1.0|0.0|RT @randyprine: Why we need Trump's tax returns. https://t.co/DUaG57942q
ujhsteacher|twitter|0.0|0.0|1.0|0.0|RT @randyprine: Why we need Trump's tax returns. https://t.co/DUaG57942q
LaOkieKat|TheTrumpLady|0.4184|0.133|0.625|0.242|"RT @TheTrumpLady: Wow! Unbelievable! #Ryan Working With Trump on Wall, Deport Criminal Illegals, Extreme Vetting, School Choice, etc. https"
DougBurges|OldeHippi|-0.7067|0.234|0.667|0.098|"RT @OldeHippi: @yashar @AndreaChalupa But, it's true!!! Nixon was nothing compared to this hell we're in right now!! Trump is a monster."
kxenp|YahBoyAhmed|0.0|0.0|1.0|0.0|RT @YahBoyAhmed: Melania Trump stole a whole speech and she on her way to becoming the First Lady but when I copy paste a paragraph on my e
madcatjo2point0|gizmodo|-0.4019|0.267|0.593|0.141|"""Donald Trump Clarifies His Plans for Destroying the Environment"" https://t.co/7j8nD2TbE5"
AnaiseRivera11|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
AnaiseRivera11|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
USATRANSEXUAL|whitebg19611|-0.5255|0.166|0.834|0.0|"RT @whitebg19611: @USATRANSEXUAL @realDonaldTrump @Maxeightyeight got to build sets, it's all Fake, it's all written, totally scripted! Tru"
sillydawg_billy|JustinRaimondo|-0.4767|0.119|0.881|0.0|"RT @JustinRaimondo: We don't need an investigation of the fake Russian ""plot"" to elect Trump: we need an investigation of the CIA spooks be"
JenJruggio|SenSanders|0.0|0.0|1.0|0.0|"RT @SenSanders: Mr. Trump may not know it, and his nominee for EPA administrator may not know it, but the debate is over. Climate change is"
lindseymfloyd|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
bonnieblue719|AriaWilsonGOP|0.4466|0.0|0.836|0.164|RT @AriaWilsonGOP: Traitors John McCain and Lindsey Graham JOIN DEMOCRATS to DELEGITIMIZE President-Elect Trump https://t.co/vqgWT8GnPr htt
bonnieblue719|truthfeed|0.4466|0.0|0.836|0.164|RT @AriaWilsonGOP: Traitors John McCain and Lindsey Graham JOIN DEMOCRATS to DELEGITIMIZE President-Elect Trump https://t.co/vqgWT8GnPr htt
HatticusFinch|twitter|-0.765|0.398|0.602|0.0|Trump is putting the country in danger. Our enemies are watching. https://t.co/jLiTCoywTw
thetinyrhino|nymag|0.0|0.0|1.0|0.0|"Just in case anyone tells you ""it's all gonna be fine."" https://t.co/1fvlSHllqe"
barney1776|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
JoinerMari|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/jWaCzABizw https://t.co/mD7GzZCYaf
JoinerMari|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/jWaCzABizw https://t.co/mD7GzZCYaf
Kitsandcrafts|youtube|-0.296|0.197|0.674|0.129|Anonymous: Trump Ability To Destroy ISIS Outlawed As Silent Coup Against Him Accelerates https://t.co/yfjsW160ly
1549321s|mcspocky|0.0|0.0|1.0|0.0|"RT @mcspocky: Liz Warren Just Made Epic Federal Move Against Trumps Corruption, Holy Sh*t [Details]  Liberal Society https://t.co/Bd11xiL"
1549321s|t|0.0|0.0|1.0|0.0|"RT @mcspocky: Liz Warren Just Made Epic Federal Move Against Trumps Corruption, Holy Sh*t [Details]  Liberal Society https://t.co/Bd11xiL"
RobertRokdawg|steph93065|-0.6636|0.243|0.757|0.0|RT @steph93065: The globalists won't give up easily. They are trying to undermine #Brexit through the courts &amp; trying to undermine Trump w/
Brooke888888|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
blueskymountain|AdamsFlaFan|-0.128|0.081|0.919|0.0|"RT @AdamsFlaFan: After Russian election rig, federal ct has precedent to install Hillary Clinton over Donald Trump https://t.co/TuSZyafGBP"
blueskymountain|dailynewsbin|-0.128|0.081|0.919|0.0|"RT @AdamsFlaFan: After Russian election rig, federal ct has precedent to install Hillary Clinton over Donald Trump https://t.co/TuSZyafGBP"
McbrideHoover|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
superdeejay64|twitter|-0.4648|0.281|0.586|0.133|"""Next eight years""How arrogant. We all know if some GOOD candidates run next election Trump is losing so hard https://t.co/kzNOA8ZCj4"
tnfortrump|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
tnfortrump|thegatewaypundit|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
loganausman|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: Durin the Army/Navy game, Trump sat on Army side in the 1st half &amp; the Navy side in the 2nd half. Obama decided to sit wi"
BurnettCynthia|LOLGOP|0.4767|0.0|0.829|0.171|RT @LOLGOP: Ways to get Trump to read intelligence briefs*Centerfolds*Highlights from Hitler speeches*Comment sections*Say they're fro
calatayud7|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
fwilson6|MarlowNYC|0.0|0.0|1.0|0.0|RT @MarlowNYC: 'Hidden Figures': The movie Trump's America needs to see https://t.co/kM3joA3g9C https://t.co/PKcgma9GFt
fwilson6|thedailybeast|0.0|0.0|1.0|0.0|RT @MarlowNYC: 'Hidden Figures': The movie Trump's America needs to see https://t.co/kM3joA3g9C https://t.co/PKcgma9GFt
grandpooba5440|datadyne007|0.431|0.0|0.875|0.125|RT @datadyne007: #SNL #WeekendUpdate perpetuating Trump's myth that CIA claimed WMDs were in Iraq. They did not. CIA was horrified Bush/Che
octaviahenke|hectormorenco|-0.6369|0.284|0.608|0.108|RT @hectormorenco: Trump should repeal and replace Obama Care for no other reason than to trash arrogant &amp; obnoxious Obama's signature dome
budnikBruce|JackDix03868724|0.5423|0.0|0.816|0.184|RT @JackDix03868724: Ex-president Vicente Fox set today Donald Trump better be careful because the food they eat is furnished by Mexico tha
wooferunleashed|MMFlint|0.0|0.0|1.0|0.0|RT @MMFlint: Trump's Sec of State: ExxonMobil CEO. That's 10 billionaires/millionaires &amp; 3 generals. Fascism's the marriage of the corp. &amp;
MoviesWorldNewz|WorldfNature|-0.6908|0.266|0.734|0.0|RT @WorldfNature: Climate Alarmist: Donald Trump Should 'Kill Himself Immediately' - Breitbart News https://t.co/ED6F9qpV4v https://t.co/XK
MoviesWorldNewz|route|-0.6908|0.266|0.734|0.0|RT @WorldfNature: Climate Alarmist: Donald Trump Should 'Kill Himself Immediately' - Breitbart News https://t.co/ED6F9qpV4v https://t.co/XK
Mhanooti|thinkprogress|0.0|0.0|1.0|0.0|RT @thinkprogress: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/uDbkj11p3M ht
Mhanooti|medium|0.0|0.0|1.0|0.0|RT @thinkprogress: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/uDbkj11p3M ht
AzizHakimiSyah|djrothkopf|0.9022|0.0|0.611|0.389|"RT @djrothkopf: Donald ""I'm, like, a smart person"" Trump ought to know that perhaps greatest sign of being smart is knowing what you don't"
johnnyb496|wagner_isabel|0.6369|0.13|0.567|0.303|"RT @wagner_isabel: New type of war? U.S. intelligence agencies have ""high confidence"" Russia acted covertly to help Trump in election https"
kleptocracynow|ezlusztig|-0.6249|0.17|0.83|0.0|"RT @ezlusztig: Purely on the basis of information publicly available - just the tip of an iceberg, presumably - Obama could devastate Trump"
SnowWhiteheart|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
SnowWhiteheart|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
INVUQT|mtracey|-0.5106|0.223|0.671|0.106|"RT @mtracey: Liberals screaming about Russia must be furious at Obama, who would've had to be complicit in the grand coverup https://t.co/Q"
INVUQT|sdrobs|-0.5106|0.223|0.671|0.106|"RT @mtracey: Liberals screaming about Russia must be furious at Obama, who would've had to be complicit in the grand coverup https://t.co/Q"
dreamyswapnil|tech2eets|0.7845|0.0|0.67|0.33|RT @tech2eets: US intelligence analysts conclude that Russia helped Trump win the 2016 elections https://t.co/x7Y992Dj90 https://t.co/Y35yt
dreamyswapnil|tech|0.7845|0.0|0.67|0.33|RT @tech2eets: US intelligence analysts conclude that Russia helped Trump win the 2016 elections https://t.co/x7Y992Dj90 https://t.co/Y35yt
RJMonstrous|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
fleshandbrand|TheBpDShow|0.0|0.0|1.0|0.0|RT @TheBpDShow: LIVE: Politics and Grits #5 | Russia Russia Russia on #spreaker #russia #trump https://t.co/0ZtRvgzQJS
fleshandbrand|spreaker|0.0|0.0|1.0|0.0|RT @TheBpDShow: LIVE: Politics and Grits #5 | Russia Russia Russia on #spreaker #russia #trump https://t.co/0ZtRvgzQJS
bulldogfinance|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
OttoBrown|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
ramrhonda|JonRiley7|-0.1531|0.143|0.738|0.119|RT @JonRiley7: Trumps Carrier deal sets a bad precedent that companies must get on Trump's good side: that's crony capitalism. https://t.c
ramrhonda||-0.1531|0.143|0.738|0.119|RT @JonRiley7: Trumps Carrier deal sets a bad precedent that companies must get on Trump's good side: that's crony capitalism. https://t.c
gailyRN|NBCPolitics|0.4019|0.0|0.803|0.197|RT @NBCPolitics: Donald Trump: I'm too smart to need daily briefings https://t.co/QXBCuXIGJF
gailyRN|nbcnews|0.4019|0.0|0.803|0.197|RT @NBCPolitics: Donald Trump: I'm too smart to need daily briefings https://t.co/QXBCuXIGJF
rockrexx|Politicringe|-0.8415|0.347|0.653|0.0|RT @Politicringe: Texas Muslim Pleads Guilty to Setting Fire to His Own Mosque (FIRST BLAMED ON TRUMP RACISM) https://t.co/0Hpg1bvv5H via @
rockrexx|breitbart|-0.8415|0.347|0.653|0.0|RT @Politicringe: Texas Muslim Pleads Guilty to Setting Fire to His Own Mosque (FIRST BLAMED ON TRUMP RACISM) https://t.co/0Hpg1bvv5H via @
AliceAl18241727|twitter|-0.1027|0.142|0.731|0.127|"Trump will give CIA  kudos when it's convenient.  When CIA might impact his election in negative way, then he berat https://t.co/s5lQVddYIh"
su_z_t|DavidYankovich|0.2732|0.0|0.909|0.091|"RT @DavidYankovich: So, Donald Trump has committed treason... This is a moment for little Marco to become Big Marco- Stand up now. https:"
MigueleSantos1|adirado29|0.6758|0.076|0.691|0.233|RT @adirado29: No one cares about the transcripts! 3 Goldman Sachs men are in Trump's Cabinet now! Does this ease your conscience at all?!
ethiojawn|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
royalviking04|Micky_Finn|-0.4019|0.13|0.87|0.0|@Micky_Finn @Kris_Sacrebleu Must be annoying to have to take off the white hood before you can sip it. https://t.co/YGyFpvTZe7
royalviking04|americannewsx|-0.4019|0.13|0.87|0.0|@Micky_Finn @Kris_Sacrebleu Must be annoying to have to take off the white hood before you can sip it. https://t.co/YGyFpvTZe7
AlwaystrumpOrg|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/JeViHG1LMG https://t.co"
AlwaystrumpOrg|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/JeViHG1LMG https://t.co"
girishglg|FoxNews|0.5423|0.0|0.774|0.226|RT @FoxNews: Trump: We're Going to Start Saying 'Merry Christmas' Again https://t.co/rFmwtKQXIZ https://t.co/PexEqzNo9E
girishglg|insider|0.5423|0.0|0.774|0.226|RT @FoxNews: Trump: We're Going to Start Saying 'Merry Christmas' Again https://t.co/rFmwtKQXIZ https://t.co/PexEqzNo9E
TommyLap77|Suntimes|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
TommyLap77|chicago|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
jrevans1963|Khanoisseur|-0.8555|0.313|0.634|0.053|"RT @Khanoisseur: Let this sink in-Trump's defense for journalists being killed in Russia:""So what, we do plenty of killing too"" https://t"
jrevans1963||-0.8555|0.313|0.634|0.053|"RT @Khanoisseur: Let this sink in-Trump's defense for journalists being killed in Russia:""So what, we do plenty of killing too"" https://t"
suzannekco|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
PrezElect_Trump|angelsofrussia|0.4359|0.0|0.869|0.131|RT @angelsofrussia: Robert is a Satan worshiper.  #robertdeniro what are you going to do now? Judge them and judge them again!!!#spiri
Mandari25733571|nytimes|-0.7096|0.258|0.742|0.0|RT @nytimes: Donald Trump ties CIA reports on Russian meddling in the election to Democrats' embarrassment over defeat https://t.co/2QMNlJ3
Mandari25733571|t|-0.7096|0.258|0.742|0.0|RT @nytimes: Donald Trump ties CIA reports on Russian meddling in the election to Democrats' embarrassment over defeat https://t.co/2QMNlJ3
Happy_Cajun|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
toilettweetage|Anomaly100|-0.5994|0.205|0.795|0.0|RT @Anomaly100: Alarm Over Witch Hunt After Trump Demands List of Civil Servants Who Worked On Climate Policy Under Obama https://t.co/KZ
toilettweetage|t|-0.5994|0.205|0.795|0.0|RT @Anomaly100: Alarm Over Witch Hunt After Trump Demands List of Civil Servants Who Worked On Climate Policy Under Obama https://t.co/KZ
cmultrading|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
TerryMcKay2|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
TerryMcKay2||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
TheGrapesOfWisc|tribelaw|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
TheGrapesOfWisc|twitter|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
Lilitree|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
RoughAcres|moderate2severe|0.0|0.0|1.0|0.0|RT @moderate2severe: #60Minutes should have asked @SpeakerRyan about Trump comparisons to Hitler. #Resist #DoYourJob Pelley! https://t.co/p
RoughAcres|paulstamatiou|0.0|0.0|1.0|0.0|RT @moderate2severe: #60Minutes should have asked @SpeakerRyan about Trump comparisons to Hitler. #Resist #DoYourJob Pelley! https://t.co/p
notthepeepspres|amma1207|0.7351|0.07|0.696|0.234|@amma1207 actions speak louder than words. What actions had trump done that proves he is a great leader? none in my book. No reason to trust
FoolishlyHigh|BernieSanders|-0.1531|0.122|0.778|0.1|RT @BernieSanders: Donald Trump is a pathological liar.  We need the help of the American people to build a movement of millions who are fo
DRHsPsychoCafe|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
DRHsPsychoCafe|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
nehadamini|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
alex_peppers|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
TOTweetFest|twitter|-0.3076|0.111|0.889|0.0|That many vote machines breaking? Why isn't this getting news attention...or did I miss it?! Part of the infrastruc https://t.co/8TXLDRaY9x
LucasGlustman|Alter_Ego_Mx|0.0|0.0|1.0|0.0|RT @Alter_Ego_Mx: #TwitterInfluence Trump on Twitter: A history of the man and his medium https://t.co/fSKJbUrWKi
LucasGlustman|linkis|0.0|0.0|1.0|0.0|RT @Alter_Ego_Mx: #TwitterInfluence Trump on Twitter: A history of the man and his medium https://t.co/fSKJbUrWKi
bheider11|billyeichner|0.6486|0.125|0.554|0.321|"RT @billyeichner: Democrats deserve better than Trump. Republicans deserve better than Trump. All Americans deserve better than this lying,"
MonicaFitz1|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
ChristineAdams3|PattiKimble|-0.6808|0.272|0.728|0.0|"RT @PattiKimble: Deride press, pull permit liberal women's group at Lincoln Memorial, enemy lists. Beginning of authoritarianismhttps://t"
randyshort|realalexjones|0.0|0.155|0.69|0.155|Megyn Kelly Blames Trump for Americans Not Trusting Mainstream Media Anymore https://t.co/ynb81jTSQk via @realalexjones
randyshort|infowars|0.0|0.155|0.69|0.155|Megyn Kelly Blames Trump for Americans Not Trusting Mainstream Media Anymore https://t.co/ynb81jTSQk via @realalexjones
jlmrbk|Stonekettle|0.4404|0.0|0.879|0.121|"RT @Stonekettle: Lately Trump supporters have taken to using the word ""cuck"" Ironically it now appears they got they themselves got cucko"
Captain_Kidd|eliasisquith|-0.7579|0.255|0.745|0.0|RT @eliasisquith: Imagine if everything Trump did during transition was intended to terrify his enemies. How would that differ from *what h
ub109ej|amjoyshow|0.0|0.0|1.0|0.0|RT @amjoyshow: .@JoyAnnReid just explained all the people linked to Donald Trump who have documented ties to #Russia and Putin #AMJoy https
NancySRed|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
MommyNooz|mommytimes|0.0|0.0|1.0|0.0|Advice to Melania Trump: Heres how to tackle cyberbullying - https://t.co/2z1IW93FNw
nakedlaughing|yashar|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
nakedlaughing|twitter|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
cherylkeats|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
MizCoretta|tonyschwartz|-0.296|0.091|0.909|0.0|RT @tonyschwartz: I don't believe anything Donald Trump says. Not one word. It is all manipulation and mind games all the time. (Same for K
SorryAbtTheFace|TheThomason|0.0|0.0|1.0|0.0|"RT @TheThomason: Realistically, I just don't know if there's time for Trump to learn to read before beginning his presidency."
realworldrj|wsj|0.4215|0.0|0.851|0.149|"This is true: Trump blasted Lockheed over out of control costs over F35s (also, not needed) https://t.co/VIV7XyGATo"
JosieRTM|kelseydarragh|-0.4404|0.176|0.758|0.066|RT @kelseydarragh: I keep acting like my problems r gunna b gone once 2016 is over but no Trump will b president and Im still gunna spend t
Dc37Deborah|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
KellsBooks|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
fahyhallowell|funder|0.0|0.0|1.0|0.0|RT @funder: Donald Trump called me David &amp; himself Goliath.I don't think he knows how that ended#TrumpIsBeingInvestigated!#TrumpLeaks
ScullyNoreen|CDZ_999|-0.8828|0.339|0.661|0.0|RT @CDZ_999: i just heard trump say he doesnt want to sit thru them . get this fuck outta contention or you are DOOMED https://t.co/3Xgk0HF
ScullyNoreen|t|-0.8828|0.339|0.661|0.0|RT @CDZ_999: i just heard trump say he doesnt want to sit thru them . get this fuck outta contention or you are DOOMED https://t.co/3Xgk0HF
Newyorker2212|Island_Canes|0.0|0.0|1.0|0.0|RT @Island_Canes: Secretary of State??? @AmbJohnBolton ... have you noticed how all these Sociopaths #trump is considering are also patholo
bebullish|nytimes|0.0|0.0|1.0|0.0|"The New Reality of TV: All Trump, All the Time, via @nytimes https://t.co/1feASpNhIG"
bebullish|nytimes|0.0|0.0|1.0|0.0|"The New Reality of TV: All Trump, All the Time, via @nytimes https://t.co/1feASpNhIG"
BlueStateBob1|mad1nola|0.0|0.0|1.0|0.0|RT @mad1nola: And why go to COMEY? Is he their go to guy for all assist for trump and his trampling of democracy! https://t.co/sJLZ7q5J5k
BlueStateBob1|twitter|0.0|0.0|1.0|0.0|RT @mad1nola: And why go to COMEY? Is he their go to guy for all assist for trump and his trampling of democracy! https://t.co/sJLZ7q5J5k
MattJSour|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
drrmittal|TuckSchool|0.0|0.0|1.0|0.0|RT @TuckSchool: Why Trump's browbeating of U.S.-based companies is a misguided approach to rebuilding jobs. https://t.co/ABo1lTmysz @Carrie
drrmittal|tuck|0.0|0.0|1.0|0.0|RT @TuckSchool: Why Trump's browbeating of U.S.-based companies is a misguided approach to rebuilding jobs. https://t.co/ABo1lTmysz @Carrie
portal4trends|twitter|-0.296|0.136|0.864|0.0|Alec Badwin levou na categoria de 'Melhor Ator Convidado' no SNL interpretando Trump. #CriticsChoice https://t.co/qcMFFykb8g
Landry777Tom|steph93065|-0.4019|0.112|0.843|0.044|"RT @steph93065: Until Jan 20, the left/MSM will do/say anything to delegitimize &amp; try to prevent Trump from taking office; their tantrum is"
going2left|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
Billandbecks|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
Billandbecks|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
HonkyTonkNights|hannity|-0.2023|0.225|0.588|0.186|WATCH: Teacher Caught On Hidden Camera Calling Trump Win An 'Act Of Terrorism' https://t.co/5lOWFzBfn9
JavyBon|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
JavyBon||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
KarmaKittySays|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
mama2fluffs|Truth247|-0.7096|0.237|0.763|0.0|RT @Truth247: Trump used 2 complain about Obama not getting intel briefings https://t.co/DhW6gAAHmS ||&amp; the arrogance will cont by him &amp; hi
mama2fluffs|huffingtonpost|-0.7096|0.237|0.763|0.0|RT @Truth247: Trump used 2 complain about Obama not getting intel briefings https://t.co/DhW6gAAHmS ||&amp; the arrogance will cont by him &amp; hi
MLorance|P0TUS|-0.3182|0.133|0.867|0.0|"RT @P0TUS: NBC News just now: ""Trump disagrees with the intel briefings that he doesn't attend"""
IlladelphAC|samsteinhp|-0.3818|0.225|0.656|0.119|@samsteinhp except when you repeat it without saying otherwise...pizza gate. You have no idea how dumb Trump supporters are
mblaber|Evan_McMullin|0.0119|0.094|0.81|0.096|RT @Evan_McMullin: It must be clear that Donald Trump is not a loyal American and we should prepare for the next four years accordingly. @r
BoringOldWhtGuy|theprospect|0.3182|0.0|0.897|0.103|"RT @theprospect: In Trump's plan, the uber-rich would see a 14% increase in after-tax income. The bottom fifth: just .07 percent. https://t"
BoringOldWhtGuy||0.3182|0.0|0.897|0.103|"RT @theprospect: In Trump's plan, the uber-rich would see a 14% increase in after-tax income. The bottom fifth: just .07 percent. https://t"
kimvie|Suntimes|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
kimvie|chicago|0.4404|0.158|0.542|0.3|"RT @Suntimes: Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
campbecc|Newyorker2212|0.3612|0.0|0.909|0.091|@Newyorker2212 He knows trump is a narcissist; he's not going to even try to stand up to him.  He's stroking his ego to make him an asset.
ciphergoth|mattyglesias|0.2617|0.057|0.786|0.157|RT @mattyglesias: Trump has a 37% approval rating. Democrats have a serious political challenge but converting Trump fans isn't it. https:/
ciphergoth||0.2617|0.057|0.786|0.157|RT @mattyglesias: Trump has a 37% approval rating. Democrats have a serious political challenge but converting Trump fans isn't it. https:/
slo220|mradamscott|0.7345|0.0|0.721|0.279|"RT @mradamscott: In short our president-elect, in cahoots with Russia, seems determined on dismantling our republic. Merry Christmas!https"
mageactivism|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
PIE20121|twitter|-0.4767|0.242|0.649|0.108|Oh Guiliani is in this to his eyeballs. He's crazy like everyone around Trump the Orange lunatic. https://t.co/SL4M5llL8N
ViterboAlberto|donfelixSPM|-0.296|0.095|0.905|0.0|"RT @donfelixSPM: Interfiri el gobierno ruso en las elecciones gringas para darle una manito a Donald Trump? l dice que no, la CIA dice q"
TimothyKopp2|Lrihendry|0.1275|0.113|0.756|0.13|RT @Lrihendry: While shopping 2day I overheard a conv with group saying isn't it great we can say Merry Christmas again &amp; not be afraid! WO
Mj4lgbtq|AJentleson|0.3472|0.0|0.904|0.096|"@AJentleson yes! It may be feel less partisan to point out Bannon, Sessions, Flynn, Pence instead of Trump, but he fits all of this!"
Mom9Ky|JoyAnnReid|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
Mom9Ky|twitter|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
buddhagirl5|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
jim_oleary|nick_dacosta|0.5859|0.0|0.648|0.352|RT @nick_dacosta: Brilliant Norwegian cartoon on #Trump https://t.co/H4amqJQCFe
jim_oleary|twitter|0.5859|0.0|0.648|0.352|RT @nick_dacosta: Brilliant Norwegian cartoon on #Trump https://t.co/H4amqJQCFe
ZappaTrustTroll|TheDemocrats|0.5514|0.0|0.818|0.182|RT @TheDemocrats: Are you:- A woman?- Under 26?Do you:- Have a pre-existing condition?- Live?- Breathe?Obamacare helps you. Don't le
cslocki|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Smallw9Victoria|KatzOnEarth|0.5106|0.0|0.852|0.148|RT @KatzOnEarth: Fun fact: The lie that Trump repeated about Obama in 2014 came from Steve Bannon's disinformation group. https://t.co/IESr
Smallw9Victoria|t|0.5106|0.0|0.852|0.148|RT @KatzOnEarth: Fun fact: The lie that Trump repeated about Obama in 2014 came from Steve Bannon's disinformation group. https://t.co/IESr
cameronhaider|apeirophobic|0.607|0.0|0.752|0.248|"@apeirophobic @NewGirl4444 that was regarding Russia's support for trump, not that Russia hacked electionPlease read next time"
JaneJanie416|POTUS|0.0986|0.248|0.421|0.331|@POTUS please save us from Trump. This is so scary
_rel8tivity_|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: Trump: 'Nobody really knows' if #ClimateChange is real. Um... Apart from every scientist who works on the subject?! Idi
RickAShepherd|youtube|0.2716|0.0|0.884|0.116|"Especially important now: Back in Sept, ABC News' Brian Ross investigated Trump's Russian, overseas business deals https://t.co/KiC6RjwGeM"
CoryKCrabtree|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
CoryKCrabtree|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
Daisypie54|DailyNewsBin|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
Daisypie54|palmerreport|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
slmbs9|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
slmbs9|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
agathawise|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
Camerannyc|NateSilver538|0.0|0.0|1.0|0.0|"RT @NateSilver538: If you're Trump, what's the rationale for picking Tillerson *other* than the Russia stuff? He's not George C. Marshall,"
FionaGillen2013|WalshFreedom|-0.6124|0.271|0.588|0.141|"@WalshFreedom Careful most of the ""people"" arguing to support Trump are Russian. Lots of fake accounts and bots out means they are worried."
caroljdavy|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
caroljdavy|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
papodedireita|chumbogrossomanaus|0.0|0.0|1.0|0.0|"Para Donald Trump reduzir as emisses de carbono prejudicam a competitividade global da Amrica e pergunta, ""Voc... https://t.co/mW24Yi9iVX"
miscelaineee|KeithOlbermann|0.0|0.0|1.0|0.0|RT @KeithOlbermann: CIA reveals how Russians ran a coup for Trump. From 10/14: the day Trump revealed he KNEW the Russians were doing it ht
WhatCandyThinks|JamesRitch1|0.656|0.0|0.856|0.144|"RT @JamesRitch1: Notice how the mood in America has changed so positively now that we know an Alpha Male is about to take charge on Jan 20,"
states37|RepublicanPunk|0.3612|0.0|0.884|0.116|"@RepublicanPunk Trump will not concede power aftee 8 years and will hold America hostage, handing power to his son, like Fidel...."
nowherenorthere|RadioFreeTom|0.0|0.0|1.0|0.0|"@RadioFreeTom If this is 'reasonable', then the 'Putin is running Trump' view can't be ruled out."
DanBoyd3|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
BrandonTozzo|davidfrum|0.296|0.0|0.872|0.128|@davidfrum so what happens if it's found Russia was helping or coordinating with the Trump campaign?
suicide_romance|elnortej|0.0|0.0|1.0|0.0|"RT @elnortej: .@SenateMajLdr kept pro-#Trump Russia hacks a secret, then Trump hired his wife, @ElaineChao. #LockHimUp #NotMyPresident"
nennaa9|YahBoyAhmed|0.0|0.0|1.0|0.0|RT @YahBoyAhmed: Melania Trump stole a whole speech and she on her way to becoming the First Lady but when I copy paste a paragraph on my e
seth_shellhouse|medium|0.0|0.0|1.0|0.0|real talk...anyone ever consider whether Donald Trump might be vilifying rural whites on purpose? #thelongcon https://t.co/IPzzStPLFi
Shanny_resqchi|MrJamesonNeat|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
Shanny_resqchi|t|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
WorldPeaceFor2|Based_Gibson|0.0|0.0|1.0|0.0|RT @Based_Gibson: TRUMP full interview at Army-Navy game https://t.co/KHlVWolzge
WorldPeaceFor2|youtube|0.0|0.0|1.0|0.0|RT @Based_Gibson: TRUMP full interview at Army-Navy game https://t.co/KHlVWolzge
maddie142519|randyprine|0.3612|0.079|0.753|0.168|"RT @randyprine: Instead of vilifying the CIA, Trump should release his taxes to prove that Russia has no incentive for helping him be elect"
BlackServative|realjunsonchan|-0.4215|0.272|0.545|0.183|RT @realjunsonchan: Brave man Joe Scarborough risks his own life to tell truth against feral idiot fake news media. #Trump #maga #underdoge
gayCAsportsfan|TomLevenson|0.0|0.0|1.0|0.0|RT @TomLevenson: It is always projection with Trump and #GOP. Always. #TrumpJunta #ClearAndPresentDanger #Resist https://t.co/zwtZlOv8D4
gayCAsportsfan|twitter|0.0|0.0|1.0|0.0|RT @TomLevenson: It is always projection with Trump and #GOP. Always. #TrumpJunta #ClearAndPresentDanger #Resist https://t.co/zwtZlOv8D4
tram03ag|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
tram03ag||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
RWNemanich|davidfrum|0.2263|0.0|0.913|0.087|"RT @davidfrum: Its true that Donald Trump doesnt have a lot of foreign policy experience, but at least hes surrounded by knowledgeable p"
GGMaury|gabrielregino|0.0|0.0|1.0|0.0|RT @gabrielregino: Y el Gabinete haciendo #RetoGuacamole y el Senado rompiendo piatas de Trump. Y la CNDH pidiendo soldados en la calle. K
AugustEve2012|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
slidewinding|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS: GOP on hill ""prepping for President Pence""-Trump investigation begins-More soon#cnn #msnbc #AMJoy #cnnsotu #this"
ScottFordTVGuy|realDonaldTrump|0.8625|0.0|0.602|0.398|"In 2017, I will respect, &amp; give @realDonaldTrump a chance. I will retract support from media &amp; talent, if they continue disrespecting Trump."
bugsy159|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
SscottSsmith84|DRUDGE_REPORT|0.2732|0.0|0.741|0.259|RT @DRUDGE_REPORT: Rick Perry Energy Secretary? https://t.co/aLPnXKPtDH
SscottSsmith84|bloomberg|0.2732|0.0|0.741|0.259|RT @DRUDGE_REPORT: Rick Perry Energy Secretary? https://t.co/aLPnXKPtDH
SerenityTau|occupydemocrats|0.4939|0.138|0.58|0.281|Dan Rather Just Called Out Fake Patriots Who Support Trumps Putin Romance In Viral Post - https://t.co/yq4LBTIkZi
MpatePat|Hotpage_News|0.3182|0.0|0.85|0.15|RT @Hotpage_News: NETANHAHU WANTS to work with #Trump on two-state solution - WASHINGTON EXAMINER https://t.co/4NbEucRxp1
MpatePat|hotpagenews|0.3182|0.0|0.85|0.15|RT @Hotpage_News: NETANHAHU WANTS to work with #Trump on two-state solution - WASHINGTON EXAMINER https://t.co/4NbEucRxp1
MsDemeanor0125|_0HOUR1|0.4588|0.0|0.769|0.231|RT @_0HOUR1: Trump should dismantle the CIA on day one :)
MaureenCKelly|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/TEGHqhLpZN https://t.co"
MaureenCKelly|thehill|0.3911|0.129|0.607|0.263|"RT @thehill: Trump suggests he doesn't need daily intelligence briefings: ""I'm, like, a smart person.""https://t.co/TEGHqhLpZN https://t.co"
elevatedgardens|yashar|0.6808|0.0|0.772|0.228|"RT @yashar: Trump's pick for Secretary of State, Exxon's Rex Tillerson, enjoying champagne toast w/ Putin + his associates after signing lu"
thenewsghetto|TurgidsonBuck|-0.7678|0.267|0.733|0.0|"@TurgidsonBuck when u say the MSM media ""fawned over Trump""- you are the one in the Twilight Zone. Even MSM doesnt agree with u lol moron"
Heidijbeck|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/qcREl7xyWa https://t.co/lZsJDdLqeo
Heidijbeck|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/qcREl7xyWa https://t.co/lZsJDdLqeo
ClaytonMuirhead|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
ClaytonMuirhead|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
MaggieMimsy|meganamram|0.0|0.0|1.0|0.0|RT @meganamram: Real question: does Trump believe in object permanence
K_DUBB_80|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
K_DUBB_80|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
AllnattChris|realDonaldTrump|-0.6478|0.249|0.751|0.0|"@realDonaldTrump @NBCNightlyNews @CNN Trump gets his intel from Putin. Trump being told to drop sanctions. Very weak, Trump."
MediaJuggernaut|ejenk|0.7906|0.0|0.696|0.304|RT @ejenk: I saw a video of Russians cheering on the rooftops in New Jersey when Trump won the election.
NonnieCon|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: Media: ""Trump's racist""""Trump's fascist""""Trump's sexist""""Trump's hitler""""Trump's a clown""""Trump's not serious"""""
B_eatrizCamargo|twitter|0.1964|0.246|0.464|0.291|Alec WON. YEEEES! Trump will be so angry! #CriticsChoice https://t.co/yUOej9hmt6
Newyorker2212|serpilcr|0.0516|0.181|0.625|0.194|"RT @serpilcr: BREAKING: Trump Attacks CIA, Defends Russia Following Intelligence Report https://t.co/RY5ZEFY77v"
Newyorker2212|reverbpress|0.0516|0.181|0.625|0.194|"RT @serpilcr: BREAKING: Trump Attacks CIA, Defends Russia Following Intelligence Report https://t.co/RY5ZEFY77v"
cosmogenesis777|worldnewsdailyreport|0.453|0.208|0.426|0.366|Now this !!!War is coming my Friend s !!!Are You ready ? https://t.co/y8F9Sraeye
Sumkindawizard|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
BladeInTheHouse|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
sabinobastidas|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
sabinobastidas|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
thisbegrm|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
ghostsirens|softbutchkate|0.9112|0.074|0.477|0.449|"RT @softbutchkate: i'm laughing bc trump is like ""his impression sucks"" yet alec won a fucking critic's choice award for it jdjdjdkdkd i lo"
rspin122112|Rex_Tillerson|0.8061|0.0|0.659|0.341|@Rex_Tillerson @ellenEspence Thank you for accepting the position! Please do right by America! Trump voters are counting on you!
mcmlynch|billmaher|-0.5859|0.266|0.592|0.141|"RT @billmaher: Its been almost a month, will I ever get used to Trump? Fuck no. Its like watching a toddler playing with a gun - you're alw"
kittens526|Vote_American|-0.1695|0.081|0.919|0.0|@Vote_American because McConnell wouldn't allow the info to be released. Now McConnell's wife has a job in Trump's cabinet. Read up
remmkm|P0TUS|-0.3182|0.133|0.867|0.0|"RT @P0TUS: NBC News just now: ""Trump disagrees with the intel briefings that he doesn't attend"""
isaacmorales559|LatestAnonNews|0.0|0.0|1.0|0.0|RT @LatestAnonNews: Meet Your New Overlordhttps://t.co/4IAynWrytn https://t.co/LnMy80BCcJ
isaacmorales559|twitter|0.0|0.0|1.0|0.0|RT @LatestAnonNews: Meet Your New Overlordhttps://t.co/4IAynWrytn https://t.co/LnMy80BCcJ
StillLes4Hill|yashar|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
StillLes4Hill|twitter|-0.5106|0.171|0.829|0.0|"RT @yashar: Carl Bernstein, of all people, saying Trump is a bigger liar than Nixon....that's something else... https://t.co/yF44LQrkI6"
gbeckyhudson|kurteichenwald|0.5574|0.0|0.847|0.153|"RT @kurteichenwald: If Trump started getting praise 4  appointments from ISIS, do you think Fox News would start running stories about how"
BroderickGreer|CBSNews|0.0|0.0|1.0|0.0|"RT @CBSNews: After seeing some of it curtailed post-Ferguson, police expect Trump to step up surplus military gear availability https://t.c"
BroderickGreer||0.0|0.0|1.0|0.0|"RT @CBSNews: After seeing some of it curtailed post-Ferguson, police expect Trump to step up surplus military gear availability https://t.c"
pinklady404|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
lorizellmill|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
codyelee|twitter|0.1786|0.0|0.918|0.082|And he doesn't have to worry about which hotel to stay at. The trump kremlin is but a whisper away. https://t.co/bSTgz0yZNb
Deteacherintell|npr|-0.1779|0.145|0.855|0.0|"As Trump Dismisses CIA, Congress Looks To Confront Russian Cyberattacks https://t.co/jYAcyr7D6W"
nightscouter|theguardian|0.0|0.0|1.0|0.0|The Republicans are delivering America into #Putin's hands. This could be our demise. #MAGA #MAGAx3 #Trumpgrets https://t.co/4Ne9UZzX2T
FMGhost09|Adenovir|-0.8658|0.386|0.614|0.0|"RT @Adenovir: Carl Bernstein, who broke the Watergate scandal that led to Nixon's resignation, said that Nixon's lies were nothing compared"
jonwasson|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
powerofpop|youtube|-0.775|0.363|0.527|0.109|Trump supporters attempting to boycott #RogueOne based on fake news. Can't make up this shit anymore. #StarWars... https://t.co/1xlDZSwEB8
Cliffor04618957|Hope012015|-0.5267|0.145|0.855|0.0|@Hope012015 @YahooNewstRump you are lying again cause I don't believe that you don't believe because you knew they were when Manafort quit
TexIrvin|SandraTXAS|-0.7906|0.389|0.611|0.0|@SandraTXAS @ReignsFreedom @skb_sara @jimlibertarian @jko417 @phil200269 @AmyMek @LodiSilverado -Terrorists that Trump will expel
JJohnson2u|ProtestDaily|-0.2263|0.119|0.881|0.0|RT @ProtestDaily: #Protest #Trump Protesters decry President-Elect Trump on International Human Rights Day - KMSP-TV https://t.co/En4rwJmVdM
JJohnson2u|fox9|-0.2263|0.119|0.881|0.0|RT @ProtestDaily: #Protest #Trump Protesters decry President-Elect Trump on International Human Rights Day - KMSP-TV https://t.co/En4rwJmVdM
MonicaFitz1|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
ledbettermark|rosierifka|0.577|0.0|0.816|0.184|"@rosierifka @PolitiFact To my knowledge, Putin does not deny the hacks, or that they were intended to favor Trump. Priebus is a null set."
JenWoodruff79|NonSnowflake|0.7506|0.0|0.632|0.368|@NonSnowflake @NutshellsGuy @trump_loves @ChastityTamu @StopStopHillary @Deneawv3Penny  Liberals love linking to Snopes. What a joke.
ktd101551|RalphHornsby|-0.4767|0.22|0.78|0.0|RT @RalphHornsby: He reads my tweets?Trump Labels CNN 'Fake News'  https://t.co/w7Doe6LNdj  #FakeNews
ktd101551|infowars|-0.4767|0.22|0.78|0.0|RT @RalphHornsby: He reads my tweets?Trump Labels CNN 'Fake News'  https://t.co/w7Doe6LNdj  #FakeNews
BitchyAmi|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
BitchyAmi|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
hgreenberg1|Left_of_Texas|-0.4215|0.229|0.706|0.065|RT @Left_of_Texas: Dan Rather: Founding Fathers warned about a demagogue president backed by a foreign adversary - https://t.co/SIQRWZL8aV
hgreenberg1|deadstate|-0.4215|0.229|0.706|0.065|RT @Left_of_Texas: Dan Rather: Founding Fathers warned about a demagogue president backed by a foreign adversary - https://t.co/SIQRWZL8aV
simi_kc88|owasow|0.128|0.104|0.769|0.127|RT @owasow: Trump claims landslide.Truth: Historic popular vote loss EC votes: 38th of 58 EC margin: 46th of 58https://t.co/jBCO
alexjonesshows|alexjonespodcast|-0.4019|0.184|0.816|0.0|Trump dismisses the CIAs claim it has evidence Russians hacked the election https://t.co/BlIQajTzOd
Moondawggie_PSN|diezesq|0.4939|0.0|0.878|0.122|RT @diezesq: My friend wants to commission anti-Trump art of Trump/Putin yaoi with Putin as the seme. Can anyone suggest an artist open for
MikeAndy128|MJB_SF|-0.6124|0.343|0.455|0.203|RT @MJB_SF: already Intelligence officials fear Trump. they need public outcry -OUR outcry - to support them. #AuditTheVote  https://t.co/5
MikeAndy128|twitter|-0.6124|0.343|0.455|0.203|RT @MJB_SF: already Intelligence officials fear Trump. they need public outcry -OUR outcry - to support them. #AuditTheVote  https://t.co/5
trulyguide|briantashman|0.128|0.118|0.739|0.143|RT @briantashman: @GoAngelo @Bencjacobs Bolton tried to blame the hacks on Bernie supporters back in July https://t.co/SdMDqRDH3b
trulyguide|mediamatters|0.128|0.118|0.739|0.143|RT @briantashman: @GoAngelo @Bencjacobs Bolton tried to blame the hacks on Bernie supporters back in July https://t.co/SdMDqRDH3b
MissLin68640163|twitter|-0.2379|0.148|0.752|0.1|"Hear, hear. Let's not just HOPE, let's work 2 guarantee there NEVER IS A tRUMP ADMINISTRATION. We R #bettertogether https://t.co/6TqVHNVPzG"
WUGolfer3118|ericgarland|-0.529|0.189|0.811|0.0|RT @ericgarland: The Russians didn't create Trump - only New York City and American gullibility could have done that.But they've got a SW
AntonioCMYK|NPR|0.1027|0.14|0.699|0.161|RT @NPR: Trump Says He Won't Sell His Businesses To Address Conflicts Of Interest https://t.co/zglt6GtTbX
AntonioCMYK|npr|0.1027|0.14|0.699|0.161|RT @NPR: Trump Says He Won't Sell His Businesses To Address Conflicts Of Interest https://t.co/zglt6GtTbX
raclibby|JoeNBC|-0.5267|0.139|0.861|0.0|@JoeNBC @maureendowd I teach my kids to take responsibility for their own behavior. Trump is here and now and lying through his teeth.
venrala|TheDemocrats|0.4939|0.0|0.802|0.198|RT @TheDemocrats: Trump has named: Anti-worker Labor SecretaryAnti-environment EPA admin.Anti-health care HHS SecretaryAnti-justice Att
DebbieW36246900|JuddLegum|-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
DebbieW36246900||-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
finbarvano|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
finbarvano||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
AminaBertarelli|mmpadellan|0.1177|0.107|0.765|0.129|RT @mmpadellan: It's not about Trump.It's not about GOP vs DEM.It's abt Nat'l Security. DEMAND investigation of #RussianHackers!https://
AminaBertarelli||0.1177|0.107|0.765|0.129|RT @mmpadellan: It's not about Trump.It's not about GOP vs DEM.It's abt Nat'l Security. DEMAND investigation of #RussianHackers!https://
calatayud7|MichaelGaree|-0.5267|0.204|0.739|0.057|"RT @MichaelGaree: Something comrade Trump's inner circle might want to consider: If he's charged with treason, guess who becomes co-conspir"
grandpooba5440|TeaPainUSA|0.128|0.092|0.797|0.112|"RT @TeaPainUSA: Trump claims the CIA said Saddam had WMDs.  Ironically, he's thinkin' of the last President that lost the popular vote."
AsapKrusty|BIackPplVines|-0.0772|0.075|0.925|0.0|RT @BIackPplVines: When Trump says he's gonna build a wall but you have a trick up your sleeve https://t.co/0kd5Bd3EO6
AsapKrusty|vine|-0.0772|0.075|0.925|0.0|RT @BIackPplVines: When Trump says he's gonna build a wall but you have a trick up your sleeve https://t.co/0kd5Bd3EO6
ChristopheJudek|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
far1762|markmobility|-0.3612|0.135|0.865|0.0|RT @markmobility: NYT Editorial: On Trump's refusal to investigate Russia. The election was indeed rigged. https://t.co/aRKMthkimV https://
far1762|nytimes|-0.3612|0.135|0.865|0.0|RT @markmobility: NYT Editorial: On Trump's refusal to investigate Russia. The election was indeed rigged. https://t.co/aRKMthkimV https://
JacquelinSusann|hectormorenco)Trump|0.25|0.113|0.722|0.165|Retweeted Hector Morenco (@hectormorenco):Trump should repeal and replace Obama Care for no other reason than... https://t.co/DqPTEb5L4L
JacquelinSusann|facebook|0.25|0.113|0.722|0.165|Retweeted Hector Morenco (@hectormorenco):Trump should repeal and replace Obama Care for no other reason than... https://t.co/DqPTEb5L4L
uniquerebel86|trump_first|-0.7845|0.299|0.56|0.141|"@trump_first He knows he has no chance  .. Murderers &amp; child molester's get plea deals all the time . heck, you can rape a child &amp; be free"
sjq11310|TearsInHeaven09|-0.5319|0.168|0.832|0.0|RT @TearsInHeaven09: LESSON:WHEN TRUMP TWEETS SOMETHING STUPIDHE IS TRYING TO MAKE YOU FORGETRUSSIA HACKED THE ELECTION FOR HIM
ABP81|michaelianblack|0.1531|0.0|0.862|0.138|@michaelianblack Bolton wishes there was evidence of Trump in his moustache
yanachoen|theatlantic|0.1027|0.224|0.517|0.259|Donald Trump's conflicts of interest: a crib sheet https://t.co/CZg1chWwAL
petabites|LBTheDemocrat|0.3367|0.0|0.888|0.112|RT @LBTheDemocrat: Obama must declassify everything the CIA has about the Russian interference before Trump is sworn in. Very important!
Smallgovtarian|ejenk|0.7906|0.0|0.696|0.304|RT @ejenk: I saw a video of Russians cheering on the rooftops in New Jersey when Trump won the election.
DebbiebB15|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
Bayathread|HappyFeminist|0.5859|0.0|0.703|0.297|@HappyFeminist follow @RachelleHodgs for brilliant graphing of Trump word salads.
t_pointe|spenser_clark|0.1017|0.122|0.667|0.211|RT @spenser_clark: Everyone is surprised that Trump is doing/saying dumb things like we didn't try to warn y'all's dumbasses over the past
AnnaHarffey|amjoyshow|-0.4404|0.132|0.868|0.0|"RT @amjoyshow: Scott Dworkin (@FUNDER) started #TrumpLeaks documenting hundreds of Trump's Russian ties, which the #FBI has denied or not r"
KlaasPeder|FoxNews..please|0.0|0.0|1.0|0.0|.@FoxNews..please wake up Mr. Trump before it is too late..
redhouse41|TheDailyEdge|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
redhouse41|twitter|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
DKWilson56|Niborobin55|-0.4416|0.154|0.846|0.0|RT @Niborobin55: @KellyannePolls @realDonaldTrump @andrewrcamp There is absolutely nothing exciting about Trump's agenda at all except his
joh53293471|jmsexton_|-0.0772|0.08|0.92|0.0|RT @jmsexton_: Three Decades Of Trump's Russian Ties Exposed In One Democratic Coalition Report https://t.co/l1MyWx1PK7 ~ @HuffingtonPost
joh53293471|huffingtonpost|-0.0772|0.08|0.92|0.0|RT @jmsexton_: Three Decades Of Trump's Russian Ties Exposed In One Democratic Coalition Report https://t.co/l1MyWx1PK7 ~ @HuffingtonPost
Hindu_League|Chellaney|-0.5106|0.121|0.879|0.0|RT @Chellaney: CIA failed to anticipate every major global event in the past 30 years. Now FBI contests its claim Russia aided Trump by hac
MattPerry1458|harrisonjp223|-0.802|0.3|0.625|0.075|RT @harrisonjp223: I hate how people are saying that star wars is anti trump just because rogue one has a female lead role. This country ha
bates_destinyy|TrillxLove|0.1531|0.088|0.802|0.111|RT @TrillxLove: RT this if trump becoming president is a nightmare and you officially lost all hope for this country. I just wanna see some
chelvis_bassman|RadioFreeTom|0.4767|0.0|0.876|0.124|"RT @RadioFreeTom: If HRC chose a SecState who ran an oil giant and got a medal from Putin, the GOPers defending Trump would re-convene the"
VaughnMKC|davebernstein|-0.2808|0.151|0.746|0.104|"RT @davebernstein: BREAKING: Donald Trump, Mitch McConnell and James Comey Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) http"
allison_lee21|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/U1KFDsn1Mf https://t.co/Z21lnE9BwB
allison_lee21|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/U1KFDsn1Mf https://t.co/Z21lnE9BwB
HeyJude_007|thenation|0.2023|0.165|0.631|0.204|RT @thenation: Donald Trump Is the Greatest Threat to American Democracy in Our Lifetime https://t.co/UJbSiEspTX
HeyJude_007|thenation|0.2023|0.165|0.631|0.204|RT @thenation: Donald Trump Is the Greatest Threat to American Democracy in Our Lifetime https://t.co/UJbSiEspTX
SaraKimbell|bostonglobe|0.0|0.0|1.0|0.0|https://t.co/XyARKcoJGs
CHURCHLADY320|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/qcREl7xyWa https://t.co/lZsJDdLqeo
CHURCHLADY320|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/qcREl7xyWa https://t.co/lZsJDdLqeo
Jodyjtaylor|Serpentine202|-0.3125|0.125|0.875|0.0|@Serpentine202 @cherrivarisco @esquire Don't be silly. He could have used the might of the USA to stop it. Or what would you have Trump do?
twistedparent|HamiltonElector|0.2298|0.123|0.757|0.12|"RT @HamiltonElector: Mr. Trump you are hardly a genius, no matter what Comrade Putin says.  We are smarter than you. We are #hamiltonelecto"
DenzildeanNY|swin24|-0.0572|0.055|0.945|0.0|"RT @swin24: Today, Trump says he doesnt want anyone hacking the U.S.In July, he called on Russia to hack the U.S. govt.https://t.co/"
RosalesRosina|losivad|-0.1779|0.209|0.606|0.185|"RT @losivad: @Nordstrom Drop all merchandise from Ivanka Trump &amp; Donald Trump, who promote racism, misogyny. Not a good look for you  #Grab"
suzannecheriton|jicastillo|-0.3818|0.148|0.852|0.0|RT @jicastillo: .@teenvogue has more balls than nearly every other news outlet covering Trump. Embarrassing. https://t.co/UVipBYrmb6
suzannecheriton|twitter|-0.3818|0.148|0.852|0.0|RT @jicastillo: .@teenvogue has more balls than nearly every other news outlet covering Trump. Embarrassing. https://t.co/UVipBYrmb6
LuciusCoverdale|misscherryjones|0.0|0.0|1.0|0.0|"RT @misscherryjones: Just when I think the CIA-Russia-Trump takes can't get any hotter, along comes John Bolton with a torch."
GrutMarge|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
CindyDcmurphy|mikandynothem|-0.5096|0.163|0.837|0.0|"RT @mikandynothem: As I drive by Trump Tower in Vegas every day, I can't help but smile. I'm reminded of the greatness America is about to"
Donna_DHKBB|SheWhoVotes|0.0|0.0|1.0|0.0|"RT @SheWhoVotes: If the Trump campaign isn't paying Paul Manafort, who is? Do you buy for 1 second he's working pro bono? #PutinTrump https"
tonic516|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: US Senators letter to Senate leaders-investigate Trump for Russian espionage#cnn #msnbc #AMJoy #cnnsotu #thiswee
revbrown51|SheriffClarke|0.0|0.0|1.0|0.0|@SheriffClarke @nytimes @washingtonpost @CNN @MSNBC @politico @HuffingtonPost Sheriff Clarke why did Trump pass you up for HLS?
SXMProgress|FwdThinking127|0.4754|0.0|0.838|0.162|"RT @FwdThinking127: Commander-in-tweet #Trump must realize he has the most powerful thumbs in the world, says @richardlevick"
Denicebrown2000|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
mms5048|SabrinaPruett|-0.2263|0.091|0.909|0.0|"RT @SabrinaPruett: @RobotSkeleton69 @Jennyrileyb @Slate The only thing Trump has is PMS, whining over news reports on Twitter. Teenagers sh"
debesponomi|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
PaulHartNYC|MMFlint|0.8689|0.077|0.568|0.355|RT @MMFlint: The CIA has determined Russia hacked into our election to help elect Donald J. Trump. Now Trump names Putin best friend as OUR
busdog|AlpertLoveday|0.0|0.0|1.0|0.0|RT @AlpertLoveday: Russian's (confirmed) involvement in our election and the personal ties to numerous members of Trump's cabinet should sc
smiley1085|vickiebd|0.0|0.0|1.0|0.0|@vickiebd @glassceiling02 @OfficialNMP Bye Trump troll
joliebeyonce|blackthought|-0.1531|0.094|0.833|0.072|"RT @blackthought: Those who are still trying to convince Trump voters he lied, what are you trying to get out of it? Real question. #sameth"
VeeVee|DRUDGE_REPORT|0.0|0.0|1.0|0.0|@DRUDGE_REPORT isn't he one of the people trump is looking to appoint? Of course he would say that.
Amertunesucre|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
Victor_bigd|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
kirmccumber|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
kirmccumber|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
xtinechau|ActionTime|0.6124|0.0|0.783|0.217|RT @ActionTime: Please Retweet:Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump #Resistance https:/
xtinechau||0.6124|0.0|0.783|0.217|RT @ActionTime: Please Retweet:Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump #Resistance https:/
LRBitisnot|dispowo|0.0|0.0|1.0|0.0|RT @dispowo: @LRBitisnot @The_Trump_Train yet he'll collect fat money for the apprentice from NBC. Hypocrisy again.NBC today show always fr
nubah2turnt|muftidank|0.7351|0.093|0.621|0.286|RT @muftidank: makeup enthusiasts must be super jealous of Trump because of how good his concealer is in covering up the word  on his f
jadeddiaspora|jazzhandmcfeels|0.1426|0.135|0.675|0.19|RT @jazzhandmcfeels: The facts: Wikileaks/DNC hacks were not Russia. RNC was not hacked by anyone. Vote fraud has been favorable to Hillary
MickBlair54|breitbart|0.128|0.0|0.857|0.143|Exclusive: Army-Navy Game Appearance 'First Day of Trump's Presidency' https://t.co/u7SL0Q9R9n
jenbrunelle2|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
AaronSMartin|sharpasahawke|0.5994|0.101|0.603|0.296|"RT @sharpasahawke: Ivanka Trump dances alone to ""Rich Girl"" by Hall and Oates, for sure."
BipsBario|nytimesworld|0.3182|0.0|0.881|0.119|RT @nytimesworld: Jerusalem mayor optimistic that Trump will relocate U.S. Embassy from Tel Aviv to Jerusalem. https://t.co/J3494K4isY http
BipsBario|nytimes|0.3182|0.0|0.881|0.119|RT @nytimesworld: Jerusalem mayor optimistic that Trump will relocate U.S. Embassy from Tel Aviv to Jerusalem. https://t.co/J3494K4isY http
shadylady1031|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
CathyNanMarie|Khanoisseur|-0.4588|0.15|0.85|0.0|RT @Khanoisseur: 2 reasons for trump rejecting daily intel briefings:1. Plausible deniability2. Busy making side deal$$ for himself @mrp
giso6150|rstevens|0.3818|0.105|0.673|0.222|"RT @rstevens: Hate to admit it, but I support Trumps choice of Cigarette Smoking Man for Surgeon General https://t.co/QDvLTsca85"
giso6150|twitter|0.3818|0.105|0.673|0.222|"RT @rstevens: Hate to admit it, but I support Trumps choice of Cigarette Smoking Man for Surgeon General https://t.co/QDvLTsca85"
K_DUBB_80|thegatewaypundit|0.6874|0.0|0.261|0.739|https://t.co/kUNwgfIJqd WELL WELL WELL..... 
Chambord22|MrDane1982|0.0|0.0|1.0|0.0|"RT @MrDane1982: The Russians were in involved assisting Bernie Sanders and Donald Trump, and now those same two are completely quite about"
rafat777|CarlaChamorros|0.0|0.0|1.0|0.0|"RT @CarlaChamorros: Vintage Trump, listen and understand why HE/WE WON:Exclusive: Donald Trump on Cabinet picks, transition process https"
ggbootsrock|meridithmcgraw|0.0|0.0|1.0|0.0|"RT @meridithmcgraw: ""I will say Donald Trump got 70 percent in Eastern Kentucky and I don't think it had anything to do with the Russians."""
PhilipAustin41|NewYorker|0.2263|0.109|0.727|0.164|RT @NewYorker: .@BorowitzReport: Poll: Americans Favor Keeping Air Force One and Cancelling Trump https://t.co/MGQdWsegjM
PhilipAustin41|newyorker|0.2263|0.109|0.727|0.164|RT @NewYorker: .@BorowitzReport: Poll: Americans Favor Keeping Air Force One and Cancelling Trump https://t.co/MGQdWsegjM
Bay_St_Wiseguy|vivelafra|-0.8977|0.373|0.627|0.0|"RT @vivelafra: This is very sinister.  What this man is describing is an Electoral College coup to unseat #Trump, no doubt exploited by #Hi"
Andy_J_Crawford|HuffPostPol|0.0|0.0|1.0|0.0|"RT @HuffPostPol: Trump says ""nobody really knows"" if climate change is real (It is.) https://t.co/zstqb4f01i https://t.co/nQg5iMdLXx"
Andy_J_Crawford|m|0.0|0.0|1.0|0.0|"RT @HuffPostPol: Trump says ""nobody really knows"" if climate change is real (It is.) https://t.co/zstqb4f01i https://t.co/nQg5iMdLXx"
I_Voted_Trump|Kentucky_Col|0.0|0.0|1.0|0.0|@Kentucky_Col 
M_F_Dupree|meganamram|0.0|0.0|1.0|0.0|RT @meganamram: Real question: does Trump believe in object permanence
bugsy159|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
slidewinding|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Letter from 17 House Dems Requesting Trump investigation#cnn #msnbc #AMJoy #cnnsotu #thisweek #resist https://t.
slidewinding||0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Letter from 17 House Dems Requesting Trump investigation#cnn #msnbc #AMJoy #cnnsotu #thisweek #resist https://t.
BurnettCynthia|downwithtyranny|0.4939|0.0|0.819|0.181|RT @downwithtyranny: Trump may name Rick Perry Energy Secretary. Perry's #1 donor: Kelcy Warren of Energy Transfer Partners-- $6 million (+
LadyTbirdRN|abbydphillip|-0.3724|0.118|0.882|0.0|"RT @abbydphillip: Trump on Fox News Sunday says he doesn't need daily intelligence briefings as POTUS because he's ""smart"" https://t.co/OUi"
LadyTbirdRN|t|-0.3724|0.118|0.882|0.0|"RT @abbydphillip: Trump on Fox News Sunday says he doesn't need daily intelligence briefings as POTUS because he's ""smart"" https://t.co/OUi"
carolefeuerman|MarkRuffalo|0.4767|0.0|0.823|0.177|"RT @MarkRuffalo: Why does Putin want Trump Pres? $500 billion opportunity for Exxon, Russia in Trump cabinet pick | MSNBC #ExxonKnew  https"
loudathelurker|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
Camplevi|FoxNews|0.4215|0.0|0.833|0.167|RT @FoxNews: Israel's Netanyahu hopes to work with Trump to undo Iran nuclear deal https://t.co/j3vPrJm5Kx
Camplevi|foxnews|0.4215|0.0|0.833|0.167|RT @FoxNews: Israel's Netanyahu hopes to work with Trump to undo Iran nuclear deal https://t.co/j3vPrJm5Kx
NetCatNews|twitter|0.0|0.0|1.0|0.0|#news #summary:  #teacher to  #trumps  #education  #pick: lets  #address the  #elephant in the  #room. its y https://t.co/36fp30p4ik
pearlohio|The_Trump_Train|-0.7783|0.694|0.306|0.0|@The_Trump_Train hell no I won't retweet
Tekki4415|politico|-0.3612|0.185|0.815|0.0|Intel world struggles to crack the code of an untrusting Trump https://t.co/sS5Y9KFskN
2tuff15|Hedge_Shot|0.5859|0.0|0.817|0.183|RT @Hedge_Shot: Bernie's Campaign Manager Shuts Down David Brock's Scapegoating of Millennials For Trump's Win via @HumanistReport https://
2tuff15||0.5859|0.0|0.817|0.183|RT @Hedge_Shot: Bernie's Campaign Manager Shuts Down David Brock's Scapegoating of Millennials For Trump's Win via @HumanistReport https://
dennis1160|FoxNews|0.0|0.0|1.0|0.0|@FoxNews Pres. Obama Hillary Russia's thing is just a way to under mind Pres. Elect Trump! America fed up with BS politics!
KeepAmerGr8|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
KellsBooks|Bluegirl_3|-0.7579|0.347|0.653|0.0|RT @Bluegirl_3: Teen Vogue editor pulls fire alarm on Trump gaslighting: He spun accusations of his falsehoods as bias https://t.co/czsi5
KellsBooks|t|-0.7579|0.347|0.653|0.0|RT @Bluegirl_3: Teen Vogue editor pulls fire alarm on Trump gaslighting: He spun accusations of his falsehoods as bias https://t.co/czsi5
dwboden|NoNo2GOP|0.34|0.106|0.721|0.173|RT @NoNo2GOP: U.S. Senate: No confirmations for Trump nominees until Obama's nominee confirmed to Supreme Court. https://t.co/7j7QmSMPGz
dwboden|change|0.34|0.106|0.721|0.173|RT @NoNo2GOP: U.S. Senate: No confirmations for Trump nominees until Obama's nominee confirmed to Supreme Court. https://t.co/7j7QmSMPGz
JHSaunders|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Uncovered-Before Donald Trump Made A Deal With Carrier, He Sued It@JoyAnnReid #obama #msnbc #cnn #dnc https://t.c"
JHSaunders||0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Uncovered-Before Donald Trump Made A Deal With Carrier, He Sued It@JoyAnnReid #obama #msnbc #cnn #dnc https://t.c"
equiibenji|ajplus|0.7778|0.0|0.746|0.254|"RT @ajplus: On January 20, 2017, Donald Trump will inherit the most sophisticated surveillance state the world has ever seen. Thanks Obama."
Chuckw12|Serpentine202|-0.1531|0.101|0.826|0.073|RT @Serpentine202: i suspect trump is barely computer-literate.but he did invite the russians to hack (not that they weren't already) http
Kat2701|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Subudhi1|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
Subudhi1|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
k_r_eckert|JuddLegum|0.34|0.0|0.906|0.094|RT @JuddLegum: 6. The American people must have the FULL STORY on Russia's role in the election before any of Trump's nat'l security nomine
bananadannas|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
JanePowers1|portersure|0.0|0.0|1.0|0.0|RT @portersure: @DaleMartin70 @Evan_McMullin @ElliottRHams it appears that foreign policy will be a business project for #trump.  it's call
jitzkow52|colinjones|-0.6048|0.225|0.775|0.0|"RT @colinjones: ""No president, including Richard Nixon, has been so ignorant of fact"" - Carl Bernstein on Trump https://t.co/5n9Z1nYRN0 htt"
jitzkow52|thedailybeast|-0.6048|0.225|0.775|0.0|"RT @colinjones: ""No president, including Richard Nixon, has been so ignorant of fact"" - Carl Bernstein on Trump https://t.co/5n9Z1nYRN0 htt"
susanwaldrop3|HamiltonElector|0.2298|0.123|0.757|0.12|"RT @HamiltonElector: Mr. Trump you are hardly a genius, no matter what Comrade Putin says.  We are smarter than you. We are #hamiltonelecto"
GustavoOrozcoH|rpp|0.0|0.0|1.0|0.0|APRENDE OE PPK!!!  Para presidir un pas hay que tener bolognas!!!   https://t.co/ofWKcqvKUD
LizKennedy_|igorvolsky|0.7003|0.0|0.775|0.225|RT @igorvolsky: I think this is exactly right and those of us resisting Trump better figure out how to effectively counter these positions.
JadeLeeea|meganamram|0.0|0.0|1.0|0.0|RT @meganamram: Real question: does Trump believe in object permanence
modurham|twitter|0.765|0.0|0.476|0.524|12 lol trump train for the win https://t.co/5MHuNpeoOe
Sabiha19Ahmed|TheDemocrats|0.505|0.0|0.824|0.176|RT @TheDemocrats: Don't forget that Donald Trump's nominee for HHS Secretary wants to repeal the law that helps millions of Americans acces
LltQuincy|ezlusztig|0.7184|0.0|0.5|0.5|RT @ezlusztig: Good thing we're friends again. https://t.co/18qMhfBGUP
LltQuincy|independent|0.7184|0.0|0.5|0.5|RT @ezlusztig: Good thing we're friends again. https://t.co/18qMhfBGUP
wasilalitaha|twitter|0.7506|0.0|0.684|0.316|Now that he won the elections Trump is now focused on things that matter to the American people https://t.co/MmhCowqOQa
softballscifi|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Scientists uncover Donald Trumps secret computer server for coordinating with the Russians https://t.co/UU7NH1fQNE via @dai
softballscifi|dailynewsbin|0.0|0.0|1.0|0.0|RT @starfirst: Scientists uncover Donald Trumps secret computer server for coordinating with the Russians https://t.co/UU7NH1fQNE via @dai
FashionHitList|ELLEmagazine|-0.8591|0.388|0.612|0.0|RT @ELLEmagazine: Teenage Girl Was Harassed and Threatened Online After Donald Trump Attacked Her on Twitter https://t.co/MBsLIAZNLi https:
FashionHitList|elle|-0.8591|0.388|0.612|0.0|RT @ELLEmagazine: Teenage Girl Was Harassed and Threatened Online After Donald Trump Attacked Her on Twitter https://t.co/MBsLIAZNLi https:
JacquelinSusann|hectormorenco|-0.6369|0.284|0.608|0.108|RT @hectormorenco: Trump should repeal and replace Obama Care for no other reason than to trash arrogant &amp; obnoxious Obama's signature dome
DiChristine|Will_Bunch|-0.7149|0.239|0.761|0.0|"RT @Will_Bunch: Worse than Watergate? Russia hacking is massive cloud over Trump presidency, and America. What caused this big mess? https:"
snarkyRedhd|twitter|0.4767|0.0|0.86|0.14|Trump - I don't have time for intelligence briefings Trump - I do have time to watch NBC news because I'm a TV new https://t.co/1BJM85GBOf
DivaDollar|NBCNews|0.4939|0.0|0.849|0.151|RT @NBCNews: Trump's cabinet picks have a combined wealth of $14.5B. How did they all make their money? https://t.co/FnfFnPNVaw https://t.c
DivaDollar|nbcnews|0.4939|0.0|0.849|0.151|RT @NBCNews: Trump's cabinet picks have a combined wealth of $14.5B. How did they all make their money? https://t.co/FnfFnPNVaw https://t.c
jjoel158|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
conservogirl|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
ARDALJONES|twitter|0.2037|0.107|0.733|0.16|Don't worry. Every few gloomy future/whiny/Trump/oil spill/extinction/moaning tweets I post a picture of a kitty. https://t.co/1xPQTtjY3q
reefwalker8|ross_marks|-0.3182|0.119|0.881|0.0|RT @ross_marks: @TheAtlantic So how many American jobs will be lost if Trump reverses the Obama-Iran nuclear deal?
kingtynk|BenghaziFour|-0.5574|0.159|0.841|0.0|RT @BenghaziFour: Obama fired General Mattis because he asked questions about Iran deal.Trump hired Mattis for the same reason. #maddog
Sbecher|DLin71|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
Sbecher|twitter|0.0|0.0|1.0|0.0|RT @DLin71: Transcript of Trump introducing John Bolton https://t.co/bO2qzG8o2k
spruceite|RubenBolling|0.0|0.0|1.0|0.0|RT @RubenBolling: Do the reasons Alexander Hamilton gave for electors to override the vote apply to Trump? Groove along to School Time Rock
DJItsMyGift|realDonaldTrump|-0.8807|0.421|0.579|0.0|@realDonaldTrump Too bad you'll be continuing your relationship with such a shitty network. Just another terrible Trump-related company.
addykateglen|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
nashvillez|McClatchyDC|0.5859|0.0|0.826|0.174|"RT @McClatchyDC: Since his election win, Trump has talked to Putin more than any other world leader https://t.co/mLBJ0589N3 https://t.co/QN"
nashvillez|mcclatchydc|0.5859|0.0|0.826|0.174|"RT @McClatchyDC: Since his election win, Trump has talked to Putin more than any other world leader https://t.co/mLBJ0589N3 https://t.co/QN"
ianabailey|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
KanwalRaja12|LethalShaam|0.5859|0.0|0.826|0.174|RT @LethalShaam: When you had enough of Russian involvement in Trump's win and you dont have the answer https://t.co/zatp4Mz90m
KanwalRaja12|twitter|0.5859|0.0|0.826|0.174|RT @LethalShaam: When you had enough of Russian involvement in Trump's win and you dont have the answer https://t.co/zatp4Mz90m
Ron_Goad|miss_adamsonn|-0.4939|0.122|0.878|0.0|@miss_adamsonn you have not provided facts that connects trump to Russia yet.  So step it up prove it.  Your blaming trump make yoyr case
DebbiebB15|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
Amertunesucre|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
ProAssad|TheEconomist|0.34|0.119|0.693|0.188|"RT @TheEconomist: Republicans are denying that Russias authoritarian, anti-American government wanted Mr Trump to win https://t.co/WGgzEMk"
ProAssad|t|0.34|0.119|0.693|0.188|"RT @TheEconomist: Republicans are denying that Russias authoritarian, anti-American government wanted Mr Trump to win https://t.co/WGgzEMk"
EFrazier512|Lrihendry|0.1275|0.113|0.756|0.13|RT @Lrihendry: While shopping 2day I overheard a conv with group saying isn't it great we can say Merry Christmas again &amp; not be afraid! WO
katlivezey|DBloom451|0.4559|0.126|0.677|0.197|RT @DBloom451: GLORIOUS DAY! Trump scored a twofer with Rex Tillerson pick as SoS: Both Liberals and @SenJohnMcCain are FREAKING OUT! Ad
meganlabrecque|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
meganlabrecque|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
kaymissman|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
kaymissman||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
angelnphx|MichaelGaree|0.0588|0.104|0.782|0.114|"RT @MichaelGaree: File under ""Don't get mad, get even."" Remember how Trump humiliated Sen. McCain? Now McCain's Senate Comm. investigating"
0ryuge|murph7041|-0.2185|0.346|0.389|0.265|"@murph7041 @RobotShlomo @jahimes @cliffschecter No Senators have alleged Trump committed treason, ya fool. :-D"
Nadia7Blue|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
robkuis|BernieSanders|-0.1531|0.122|0.778|0.1|RT @BernieSanders: Donald Trump is a pathological liar.  We need the help of the American people to build a movement of millions who are fo
tonic516|FreddyLawrence1|-0.0772|0.105|0.801|0.094|"RT @FreddyLawrence1: This is spot on.It's up to @POTUS if he wants a legacy, or to have Trump finish him off being disgraced w:own party di"
RamblingDon|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
LauraStevensWSJ|rebeccaballhaus|0.2263|0.0|0.888|0.112|RT @rebeccaballhaus: Trump admin picks so far:- 3 billionaires- 5 millionairesTotal net worth: close to $10B https://t.co/ITS2uRIgpV htt
LauraStevensWSJ|wsj|0.2263|0.0|0.888|0.112|RT @rebeccaballhaus: Trump admin picks so far:- 3 billionaires- 5 millionairesTotal net worth: close to $10B https://t.co/ITS2uRIgpV htt
Rajivkapoor2318|Newsmax|-0.25|0.133|0.867|0.0|Michael Moore Plans to Protest at Trump Inauguration https://t.co/NLYMXzYmVq via @Newsmax Moore is a buffoon
Rajivkapoor2318|newsmax|-0.25|0.133|0.867|0.0|Michael Moore Plans to Protest at Trump Inauguration https://t.co/NLYMXzYmVq via @Newsmax Moore is a buffoon
MpatePat|mitchellvii|0.2732|0.0|0.851|0.149|RT @mitchellvii: Report: Rick Perry on Trump's Energy Secretary Short List - Breitbart https://t.co/zcphgxiv2n
MpatePat|breitbart|0.2732|0.0|0.851|0.149|RT @mitchellvii: Report: Rick Perry on Trump's Energy Secretary Short List - Breitbart https://t.co/zcphgxiv2n
DykesJeanie|ABC|-0.3818|0.354|0.488|0.159|@ABC @BrianRoss Hail King Trump :(
SocialTwurker|Lollardfish|0.4215|0.0|0.891|0.109|"RT @Lollardfish: ""What did you do when Trump installed his empire, grandpa?""""I used my media power to yell at liberal students to be nice"
biotrooferredux|noclador|0.0|0.0|1.0|0.0|RT @noclador: #Trump transition team meeting to discuss the next head of the @CIA... https://t.co/rbCZZjJPiC
biotrooferredux|twitter|0.0|0.0|1.0|0.0|RT @noclador: #Trump transition team meeting to discuss the next head of the @CIA... https://t.co/rbCZZjJPiC
Ocande|EccehomoSetrina|0.0|0.0|1.0|0.0|RT @EccehomoSetrina: Ya Trump escogi director de la DEA. #SNL https://t.co/eOoz1CiqH2
Ocande|twitter|0.0|0.0|1.0|0.0|RT @EccehomoSetrina: Ya Trump escogi director de la DEA. #SNL https://t.co/eOoz1CiqH2
lauowolf|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
Ben4Pres2020|Tina49747372|-0.0516|0.128|0.752|0.119|@Tina49747372 @Perpetual_Now All the smart Republicans are keeping their distance. The next Trump scandal is just around the corner.
FakeDanTosello|WalshFreedom|0.4939|0.076|0.725|0.198|"@WalshFreedom I'm glad you stuck to your principles, btw... not that my opinion matters.But yeah, Trump didn't have them to begin with."
gbeckyhudson|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
kootnikoff|thehill|0.4767|0.0|0.853|0.147|#Putin tells him all he needs to know: #Trump on intelligence briefings: 'I get it when I need it' https://t.co/egknwlyMvO
canada_panda|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
NicoleCynLane|twitter|0.0|0.0|1.0|0.0|LoL...poor Mr. Trump...can't catch a break! https://t.co/FIl5v5NyLo
LaurelSnyder|VoteHillary2016|0.0|0.0|1.0|0.0|"RT @VoteHillary2016: Trump's Secretary of State pick, @Exxon's @rex_tillerson, toasting Putin &amp; associates after signing lucrative deal. ht"
cwegan|JoeNBC|0.3612|0.0|0.889|0.111|RT @JoeNBC: The first time Donald Trump and Condi Rice spoke was when she called to recommend Rex Tillerson for State.
EclecticArts2|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
Tamaraciocci|melreynoldsU|0.5423|0.0|0.809|0.191|RT @melreynoldsU: Please retweet @HillaryClinton and urge her to say something publicly about the Russians helping Trump. We need her voice
koalaqueen53|tribelaw|-0.3612|0.111|0.889|0.0|"RT @tribelaw: This is gravely disquieting. @EllenLWeintraub is an impeccable source, and what she says about Trump's White House Counsel is"
Tull007|JuddLegum|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
Tull007|t|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
joh53293471|USARedOrchestra|0.0|0.0|1.0|0.0|"RT @USARedOrchestra: CT Rep. Jim Himes call Trump ""completely unhinged"" and calls for the electoral college to do what it was designed for."
boweryboyz|helenmaryme|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
boweryboyz|twitter|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
SicSemprSeattle|thehill|0.0|0.0|1.0|0.0|"RT @thehill: Trump, lawmakers split on severity of Russian election interferencehttps://t.co/ZUkh3Tv82j https://t.co/VcHo3HAfGQ"
SicSemprSeattle|twitter|0.0|0.0|1.0|0.0|"RT @thehill: Trump, lawmakers split on severity of Russian election interferencehttps://t.co/ZUkh3Tv82j https://t.co/VcHo3HAfGQ"
carlosdz|CNET|0.0|0.0|1.0|0.0|"RT @CNET: On SNL, 'Breaking Bad's Walter White joins Trump cabinet https://t.co/IypAGpsth1 https://t.co/NOSHn0v02S"
carlosdz|cnet|0.0|0.0|1.0|0.0|"RT @CNET: On SNL, 'Breaking Bad's Walter White joins Trump cabinet https://t.co/IypAGpsth1 https://t.co/NOSHn0v02S"
benthere536|BrianWestrate|0.4118|0.0|0.861|0.139|"@BrianWestrate Mr. Westrate, with Russian interference to elect Trump, what do you think of this? Value your input.https://t.co/2TMpDMsNKy"
venrala|sierraclub|-0.2144|0.093|0.907|0.0|"RT @sierraclub: Trump's cabinet represents a who's who of climate-deniers and fossil fuel hacks, so #Tillerson's selection is shocking, but"
shbeaty|twitter|-0.0572|0.064|0.936|0.0|Another reason why I don't want Bolton to have ANY part in Trump government.  I remember his performance under G. W https://t.co/R0ssa55BqZ
DrDejnozka|immigrant4trump|0.4404|0.081|0.769|0.15|"RT @immigrant4trump: President Trump is Going to Make America Great Again Regardless of the Color of Your Skin, No More Business As Usual G"
mammothfactory|jon_bois|0.0|0.0|1.0|0.0|"RT @jon_bois: These next four years, were going to need to oppose Donald Trump at every turn. Lets get started  now. https://t.co/pW4ekS"
mammothfactory|t|0.0|0.0|1.0|0.0|"RT @jon_bois: These next four years, were going to need to oppose Donald Trump at every turn. Lets get started  now. https://t.co/pW4ekS"
ursulasalcove|RuthHHopkins|0.5859|0.0|0.847|0.153|RT @RuthHHopkins: Russia helped Trump win. The CIA has confirmed this. The election is invalid. There's opinions &amp; there's facts. This is f
cocktailgurl17|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
cocktailgurl17||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
lindadoherty4|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
SecularLad|z0mgItsHutch|-0.765|0.223|0.777|0.0|@z0mgItsHutch If they knew Trump had plans to start a nuclear war they might lie about it. As a tech guy it's not likely they were hacked.
remmkm|paul_lander|0.1531|0.098|0.781|0.121|"RT @paul_lander: Trump is now fighting with the CIA, look for him to start new intelligence agency with Putin called the KKKGB"
susanmanners|YouTube|0.0|0.0|1.0|0.0|Weekend Update: Angela Merkel on Donald Trump - SNL https://t.co/tef78inEN8 via @YouTube  #loveAngela
susanmanners|youtube|0.0|0.0|1.0|0.0|Weekend Update: Angela Merkel on Donald Trump - SNL https://t.co/tef78inEN8 via @YouTube  #loveAngela
Sunny_Tag|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
JohnHen39949447|DanScavino|0.0|0.0|1.0|0.0|@DanScavino not going to happen under a Trump watch !
NioviEducation|MMFlint|0.0|0.0|1.0|0.0|RT @MMFlint: Trump's Sec of State: ExxonMobil CEO. That's 10 billionaires/millionaires &amp; 3 generals. Fascism's the marriage of the corp. &amp;
NeedsMore_Walt|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
slsall|thehill|0.0|0.0|1.0|0.0|RT @thehill: Trump goes after NBC news in tweethttps://t.co/32I8myfDsw https://t.co/vj13vixfUJ
slsall|twitter|0.0|0.0|1.0|0.0|RT @thehill: Trump goes after NBC news in tweethttps://t.co/32I8myfDsw https://t.co/vj13vixfUJ
Bellalindafox|smartinez411|0.1779|0.0|0.898|0.102|"RT @smartinez411: How long before Trump convinces armed trolls to ""self investigate"" NBC News #Resist https://t.co/FDoYKzOsCW"
Bellalindafox|twitter|0.1779|0.0|0.898|0.102|"RT @smartinez411: How long before Trump convinces armed trolls to ""self investigate"" NBC News #Resist https://t.co/FDoYKzOsCW"
MarisolR0515|FINALLEVEL|0.9324|0.0|0.429|0.571|"RT @FINALLEVEL: FYI: I dont Block FLTG Trump supporters They like ME, so they cant be ALL bad  lol"
Willie_Jacobsz|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
KeepAmerGr8|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
cubsb4bears|bannerite|0.5267|0.0|0.833|0.167|@bannerite @RexHuppke @DapperSuppIy @realDonaldTrump Trump will put this on and tell us stories about his courageous military experiences.
LoriWill213|therealcornett|0.0|0.0|1.0|0.0|RT @therealcornett: Drip Drip: Activist Who Served on George Soros-Financed Boards Behind Scheme to Take Trumps Electoral College Votes ht
YourDailyKarmaa|yourdailykarma|0.4215|0.0|0.797|0.203|Netanyahu hopes to work with Trump to undo Iran nucleardeal https://t.co/WoAr8yT39t https://t.co/VoG32R85wO
monahb|KFILE|0.5719|0.0|0.871|0.129|@KFILE that is so absurd that I don't understand why Politico would give it any air at all.  Ex. of why Trump won - media took bait again
xkr99|KiaraMistisses|0.3182|0.0|0.796|0.204|@KiaraMistisses @ScottPresler And I am sure Trump would say #FuckKiaraMistisses also....
YankyNussen|twitter|0.0|0.0|1.0|0.0|The headline should've read; Trump will work with Israel to eliminate Iran's nuclear system from the face of the ea https://t.co/EtWpYRfUnq
DavidKARE11|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
MBarber84211320|Jxnewton|0.1027|0.12|0.741|0.139|"RT @Jxnewton: Oh look, an Australian pol advertising Trump Hotel.No conflicts of interest here. Move on folks.@kurteichenwald @Fahrentho"
wotshaking|whatshaking|-0.5859|0.407|0.593|0.0|"Where Trump Critics See Conflicts, Partners See GoldenOpportunities https://t.co/WamHcUeVO5"
mikey_who_|twitter|0.0|0.0|1.0|0.0|By now we should have realized that the only thing that will work on the 3 year old that is Trump is reverse psycho https://t.co/HZrxbdt4fF
IbisTerry|mikandynothem|0.3802|0.088|0.767|0.146|RT @mikandynothem: Ruth Bader Ginsburg said she would resign if Trump won. Hit the road lady! That will give Trump even more Conservatives
constantino_sam|pinterest|-0.4648|0.216|0.784|0.0|Give Hillary's Dad a Condom - ANTI HILLARY PRO TRUMP POLITICAL BUMPER STICKER https://t.co/bupz1ZTsPG
zebrasnake|jojoh888|0.0|0.0|1.0|0.0|@jojoh888 @Deplorable_JJ but trump let the dogs out woof woof woof woof
piresl|AP4LP|0.3244|0.0|0.885|0.115|"RT @AP4LP: Liberal Logic: ""You dont need assault rifles. Govt wont turn tyrannical but Trump is the next Hitler!"""
rossetti_nancy|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
MJBodary|sodagrrl|-0.6597|0.221|0.779|0.0|RT @sodagrrl: Brian Williams Takes a Hypocritical Shot at Trump and Can't Get out of the Line of Fire Fast Enough https://t.co/rDbZRgHwbA
MJBodary|ijr|-0.6597|0.221|0.779|0.0|RT @sodagrrl: Brian Williams Takes a Hypocritical Shot at Trump and Can't Get out of the Line of Fire Fast Enough https://t.co/rDbZRgHwbA
cellaruve25|politicususa|0.3182|0.09|0.758|0.152|RT @politicususa: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests via @politicususa https://t.co/IKDOxKghqQ #p2 #c
cellaruve25|politicususa|0.3182|0.09|0.758|0.152|RT @politicususa: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests via @politicususa https://t.co/IKDOxKghqQ #p2 #c
odesssatweets|gwatsky|0.0|0.0|1.0|0.0|RT @gwatsky: Trump cabinet really coming together https://t.co/RxpDahvTA5
odesssatweets|twitter|0.0|0.0|1.0|0.0|RT @gwatsky: Trump cabinet really coming together https://t.co/RxpDahvTA5
srfcwaffles|FoxNews|0.0772|0.0|0.92|0.08|RT @FoxNews: GOP senators challenge Trump over secretary of state prospect's Russia ties https://t.co/UqUGC6Lvoh via @foxnewspolitics
srfcwaffles|foxnews|0.0772|0.0|0.92|0.08|RT @FoxNews: GOP senators challenge Trump over secretary of state prospect's Russia ties https://t.co/UqUGC6Lvoh via @foxnewspolitics
capitalist_king|TheStreet|-0.4522|0.165|0.835|0.0|RT @TheStreet: What gay Americans and undocumented workers really stand to lose under Trump: https://t.co/tPaifxJd0b https://t.co/XaLm9VcK4i
capitalist_king|thestreet|-0.4522|0.165|0.835|0.0|RT @TheStreet: What gay Americans and undocumented workers really stand to lose under Trump: https://t.co/tPaifxJd0b https://t.co/XaLm9VcK4i
WellsCharlene|mitchellvii|0.2732|0.0|0.851|0.149|RT @mitchellvii: Report: Rick Perry on Trump's Energy Secretary Short List - Breitbart https://t.co/zcphgxiv2n
WellsCharlene|breitbart|0.2732|0.0|0.851|0.149|RT @mitchellvii: Report: Rick Perry on Trump's Energy Secretary Short List - Breitbart https://t.co/zcphgxiv2n
dpkphdcpt|nprpolitics|0.0|0.0|1.0|0.0|RT @nprpolitics: FACT CHECK: Trump Claims A 'Massive Landslide Victory'  But History Differs https://t.co/vIRCDk4TX1
dpkphdcpt|npr|0.0|0.0|1.0|0.0|RT @nprpolitics: FACT CHECK: Trump Claims A 'Massive Landslide Victory'  But History Differs https://t.co/vIRCDk4TX1
WendyJFluga28|WayneRoot|0.3481|0.0|0.891|0.109|"RT @WayneRoot: Fed will raise rates 4 ""Trump Economy""? So they admit they've kept rates at 0 for 8 yrs because of ""Obama economy?""https://"
WendyJFluga28||0.3481|0.0|0.891|0.109|"RT @WayneRoot: Fed will raise rates 4 ""Trump Economy""? So they admit they've kept rates at 0 for 8 yrs because of ""Obama economy?""https://"
conserveguitar|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
modernbob|helenmaryme|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
modernbob|twitter|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
NylaNorris|TheDonaldNews|0.128|0.111|0.754|0.136|RT @TheDonaldNews: FBI Investigation Refutes CIA=&gt; Theres No Evidence Russia Tried to Help Trump https://t.co/lUPBb1wd0y #FoxNews #Tucker
NylaNorris|thegatewaypundit|0.128|0.111|0.754|0.136|RT @TheDonaldNews: FBI Investigation Refutes CIA=&gt; Theres No Evidence Russia Tried to Help Trump https://t.co/lUPBb1wd0y #FoxNews #Tucker
carlyle65270|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
carlyle65270|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
SusieSpirit38|HowBoutAMartini|0.0|0.0|1.0|0.0|"@HowBoutAMartini @redsteeze When you have a puppet in Trump, who wouldn't?"
MATUGAMATUGA|YourAnonCentral|-0.4939|0.144|0.856|0.0|"RT @YourAnonCentral: Steal this: Open Call for mobilization against the inauguration of Donald #Trump on January 20, 2017 #DisruptJ20  http"
girishglg|FoxNews|-0.296|0.145|0.855|0.0|"RT @FoxNews: .@ericbolling: Trump to Stop 'Banksters', CEOs From 'Fooling' Average Americans https://t.co/MvCy3Ou08b https://t.co/Mq5RkPThrV"
girishglg|insider|-0.296|0.145|0.855|0.0|"RT @FoxNews: .@ericbolling: Trump to Stop 'Banksters', CEOs From 'Fooling' Average Americans https://t.co/MvCy3Ou08b https://t.co/Mq5RkPThrV"
PalbaySpyshots|gizmodo|0.8481|0.0|0.662|0.338|And #CNN #MSNBC et al...tried to help Trump LOSE...So What? CIA Report Concludes That Russia Tried to Help Trump Win https://t.co/Ttqfr0WMeQ
waldmania|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
greggypoo65|carolinagirl63|0.5994|0.0|0.794|0.206|RT @carolinagirl63: It was beautiful to see. Army-Navy Game Appearance 'First Day of Trump's Presidency' https://t.co/hAuw7zjdbE
greggypoo65|breitbart|0.5994|0.0|0.794|0.206|RT @carolinagirl63: It was beautiful to see. Army-Navy Game Appearance 'First Day of Trump's Presidency' https://t.co/hAuw7zjdbE
danknapp76|feliciaw5853|-0.2263|0.148|0.742|0.109|"RT @feliciaw5853: Obama trapped in presidency defining moment. Like Lincoln, unavoidable decision. Have CIA release intel on Trump. https:/"
danknapp76||-0.2263|0.148|0.742|0.109|"RT @feliciaw5853: Obama trapped in presidency defining moment. Like Lincoln, unavoidable decision. Have CIA release intel on Trump. https:/"
ont2alb|TrumpNewMedia|0.4648|0.0|0.856|0.144|RT @TrumpNewMedia: IS #GEORGESOROS EVER GOING TO BE HELD RESPONSIBLE FOR HIS  #CRIMES?  #Reuters #NeverRomney #Bloomberg #NBCNews #Trump #M
dbly|stateinnovation|0.0|0.0|1.0|0.0|"RT @stateinnovation: WATCH: @nick_rathod joins @amjoyshow to discuss #NCgov and how states must organize to resist, counter #Trump https://"
dbly||0.0|0.0|1.0|0.0|"RT @stateinnovation: WATCH: @nick_rathod joins @amjoyshow to discuss #NCgov and how states must organize to resist, counter #Trump https://"
deepakkhurana|NYMag|-0.3612|0.163|0.837|0.0|RT @NYMag: New York City will continue to be itself  a theater of freaks and refugees and the restless https://t.co/6R26ySgY3d #RTLNY
deepakkhurana|nymag|-0.3612|0.163|0.837|0.0|RT @NYMag: New York City will continue to be itself  a theater of freaks and refugees and the restless https://t.co/6R26ySgY3d #RTLNY
JamesGreenBronx|ClydeHaberman|-0.296|0.091|0.909|0.0|"RT @ClydeHaberman: Trump team says he had 1 of ""biggest Electoral College victories in history."" In fact, his % of electors puts him No. 46"
1finekitty|donnabrazile|0.0|0.155|0.69|0.155|RT @donnabrazile: CIA report: Russia hacked the Democrats to help Trump https://t.co/P6nCbMMAvP via @voxdotcom
1finekitty|vox|0.0|0.155|0.69|0.155|RT @donnabrazile: CIA report: Russia hacked the Democrats to help Trump https://t.co/P6nCbMMAvP via @voxdotcom
lovesnlwomen|softbutchkate|0.9112|0.074|0.477|0.449|"RT @softbutchkate: i'm laughing bc trump is like ""his impression sucks"" yet alec won a fucking critic's choice award for it jdjdjdkdkd i lo"
rudikolenc|nytimesworld|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
rudikolenc|nytimes|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
grandpooba5440|JanaBlade1|-0.34|0.094|0.906|0.0|"RT @JanaBlade1: ""FBI and CIA"" First mistake was allowing trump to run w/out showing his tax returns. That would offer much needed info into"
SweeetSpot|KeithOlbermann|0.0|0.0|1.0|0.0|RT @KeithOlbermann: CIA revealed Russia HAD tampered for Trump. From 10/14: that time Trump revealed he knew they were doing it for him htt
bachic2|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
tampadougw|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
TheCorollary|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
TheCorollary||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
MetaphorMirror|FoxNews|0.4215|0.0|0.843|0.157|RT @FoxNews: Israel's Netanyahu hopes to work with Trump to undo Iran nuclear deal https://t.co/3YTZNxycM1 https://t.co/JGo5xpEfth
MetaphorMirror|foxnews|0.4215|0.0|0.843|0.157|RT @FoxNews: Israel's Netanyahu hopes to work with Trump to undo Iran nuclear deal https://t.co/3YTZNxycM1 https://t.co/JGo5xpEfth
bobshell1968|The_Last_NewsPa|0.6249|0.0|0.769|0.231|@The_Last_NewsPa @Snoopy_thats_me trump is coming. It will all be restored to American values. Not libtards ways of last 8 yrs
ladybuggedhc|420weedin|0.0516|0.134|0.722|0.144|RT @420weedin: Trump's attorney general pick threatens years of progress in marijuana reform #legalizeIT #marijuana https://t.co/CsUBoFfxjZ
ladybuggedhc|dailykos|0.0516|0.134|0.722|0.144|RT @420weedin: Trump's attorney general pick threatens years of progress in marijuana reform #legalizeIT #marijuana https://t.co/CsUBoFfxjZ
Manyi5|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
JHSaunders|KyleNeven1|-0.5672|0.162|0.838|0.0|RT @KyleNeven1: #trumpvoterregrets cracking me up! They r finally realizing #Putin owns #Trump. #TrumpLeaks r gonna slay this fool &amp; his fl
wendellshaw5|JasonMillerinDC|0.0|0.0|1.0|0.0|RT @JasonMillerinDC: Trump's education secretary pick plans to get rid of Common Core standards https://t.co/Xx1DYeSV8G via @nypost
wendellshaw5|nypost|0.0|0.0|1.0|0.0|RT @JasonMillerinDC: Trump's education secretary pick plans to get rid of Common Core standards https://t.co/Xx1DYeSV8G via @nypost
Ranthruredlight|jdakwar|-0.8779|0.387|0.613|0.0|"RT @jdakwar: Horrific genocidal statement by military veteran and former congressman Allen West, a notorious Muslim hater emboldened by Tru"
ridgway_kelsey|TheDemocrats|0.5514|0.0|0.818|0.182|RT @TheDemocrats: Are you:- A woman?- Under 26?Do you:- Have a pre-existing condition?- Live?- Breathe?Obamacare helps you. Don't le
pisannd5|kurteichenwald|0.7089|0.0|0.772|0.228|"RT @kurteichenwald: Trump says: So smart doesnt need daily intel briefings, knows more about ISIS than military, knows tax code better than"
RazorCabron|kayfabenews|0.0|0.0|1.0|0.0|https://t.co/JTDvqZ686P #MAGA #WWE #TNA
lIl0IlI|intlspectator|-0.3818|0.254|0.595|0.151|RT @intlspectator: 2016- Trump win- Brexit- Italy referendum fail- Syria- Turkey coup attempt- N Korea nuclear tests- ISIS attacks
SocialPowerOne1|politicususa|0.3182|0.126|0.662|0.212|Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests https://t.co/Eghd6ic7s8
Mrwilbury|benschwartzy|-0.5177|0.218|0.66|0.122|"RT @benschwartzy: It only took one FBI agent to ruin Nixon (Felt) and one to ruin Hillary (Comey). So, I'm very happy to see Trump making a"
artopb|Mr_Bukowski|0.0|0.0|1.0|0.0|"RT @Mr_Bukowski: Y gracias a Donald Trump, esta familia estar unida el da de la fiesta.https://t.co/DFQftPFVrW"
KellsBooks|MrJamesonNeat|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
KellsBooks|t|-0.4404|0.255|0.607|0.138|RT @MrJamesonNeat: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/wv
CSTearlyoften|chicago|0.4404|0.175|0.492|0.333|"Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/N9TPzxRqFI https://t.co/akKz3f6Ciw"
Suntimes|chicago|0.4404|0.175|0.492|0.333|"Lynn Sweet: Trump rejects CIA intelligence on Russia, daily briefings https://t.co/4orXTJrwfP https://t.co/hIZtjOwZNF"
wetsprocket|tomtomorrow|-0.7841|0.247|0.703|0.05|RT @tomtomorrow: Thought of what Trump's election means for this country has left me feeling the sort of grief I have felt after death of s
Steven_Strauss|justinhendrix|0.0|0.0|1.0|0.0|@justinhendrix @JuddLegum @thinkprogress I bet trump repeats this before tomorrow morning
iAbu3adel|youtube|0.0|0.0|1.0|0.0| SNL: Bryan Cranston's 'Walter White' named DEA chief in Trump's cabinet https://t.co/8AdUDDSUxO
Kylerob28|Ckzoote|-0.5423|0.132|0.868|0.0|@Ckzoote @birbigs not this chicken hawk you post about this mug in every trump thread are you selling them or something? Go fuck yourself
PeterBacon5|GoAngelo|0.5106|0.0|0.858|0.142|"RT @GoAngelo: And a few days later, he excitedly posted on his facebook page that the Trump administration will ""exterminate"" all muslims h"
MarlaJ101|BettyBowers|0.9169|0.0|0.578|0.422|"RT @BettyBowers: Trump is like a smart person in the same sense he is like a modest person, or an honest person, or a faithful person or"
PhiKapMom|RepAdamSchiff|-0.34|0.118|0.882|0.0|RT @RepAdamSchiff: There's overwhelming evidence of Russian hacking of our elections. By denying it Trump has essentially become a propagan
nancychatter|twitter|0.6759|0.0|0.754|0.246|"This is a person who doesn't know, he ""don't"" realize that stupid is as stupid does.His tweets personifies ""Trump https://t.co/PWwaxgRZDs"
oufenix|tomtomorrow|-0.3182|0.182|0.704|0.114|"RT @tomtomorrow: Trump's  victory is as if your loved one died, and you grieve, and then they are brought back to life the next day and kil"
cjthefineartist|cjthefineartist|-0.8353|0.308|0.692|0.0|"RT @cjthefineartist: Trump cannot ethically take the oath. He cannot protect us from any enemies, when he is the enemy from within #RussiaH"
otohp|AP|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
otohp|t|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
AJ_Rutten|Atul_Gawande|0.4878|0.096|0.659|0.245|"RT @Atul_Gawande: Dept of This-Isn't-SNL. Trump: I don't need daily security briefings because ""I'm, like, a smart person"" https://t.co/9N8"
AJ_Rutten|t|0.4878|0.096|0.659|0.245|"RT @Atul_Gawande: Dept of This-Isn't-SNL. Trump: I don't need daily security briefings because ""I'm, like, a smart person"" https://t.co/9N8"
bait51|absolutelyhats|-0.5267|0.134|0.866|0.0|RT @absolutelyhats: @wycats 4. Be very vocal in every forum available 2 us when we observe Trump's violations of our rights &amp; our democracy
Donna_DHKBB|SheWhoVotes|0.0|0.0|1.0|0.0|RT @SheWhoVotes: Article notes Manafort may still be on retainer for Putin's Ukraine goon; note also that Trump's not paying Manafort https
maddog301|MaxAbrahms|0.0|0.0|1.0|0.0|"RT @MaxAbrahms: Officials familiar with briefings given to Congress say CIA assessment ""wasn't as definitive as has been portrayed."" https:"
dvrjr|childoflight4|-0.6597|0.302|0.554|0.144|"RT @childoflight4: 30% of Latinos (like me) LOVE Donald Trump yet these racist race baiting liars keep claiming its ""white people"" STOP THE"
sleepyjoe2|DRUDGE_REPORTKnuckleheads|0.6369|0.086|0.591|0.323|@DRUDGE_REPORTKnuckleheads like #JohnBolton want to drag America into a fact free #Trump alternate reality where nothing is real.
plowman_robert|immigrant4trump|-0.6597|0.231|0.769|0.0|"RT @immigrant4trump: Video: CNN Goes Nuts Over Russians &amp; Fake News, hacks cites Buzzfeed as their source #Maga #Trump https://t.co/SnpTgmY"
plowman_robert|t|-0.6597|0.231|0.769|0.0|"RT @immigrant4trump: Video: CNN Goes Nuts Over Russians &amp; Fake News, hacks cites Buzzfeed as their source #Maga #Trump https://t.co/SnpTgmY"
Amsoflyy|MMFlint|0.8689|0.077|0.568|0.355|RT @MMFlint: The CIA has determined Russia hacked into our election to help elect Donald J. Trump. Now Trump names Putin best friend as OUR
slmbs9|JulieAnnLily|-0.3818|0.106|0.894|0.0|RT @JulieAnnLily: @robreiner We need emergency filing to halt EC. We have Russia interference &amp; collusion w trump &amp; trump team and GOP lead
Tull007|JuddLegum|-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
Tull007||-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
WorldwideHerald|business|-0.34|0.167|0.833|0.0|RT @business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/6l8izhUs9D https://t.co/0drSTTUrnr
WorldwideHerald|bloomberg|-0.34|0.167|0.833|0.0|RT @business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/6l8izhUs9D https://t.co/0drSTTUrnr
Andy_J_Crawford|CNNPolitics|0.0|0.0|1.0|0.0|"RT @CNNPolitics: Donald Trump: ""Nobody really knows"" if climate change is real https://t.co/BQ4z69MJJn https://t.co/Z9xI0BZ4Jt"
Andy_J_Crawford|cnn|0.0|0.0|1.0|0.0|"RT @CNNPolitics: Donald Trump: ""Nobody really knows"" if climate change is real https://t.co/BQ4z69MJJn https://t.co/Z9xI0BZ4Jt"
NedSparks|Psyllius|-0.5267|0.236|0.764|0.0|@Psyllius They worked together. You are lying if you say they didn't.https://t.co/cmrMwPlkql
democrat_mn|HamiltonElector|-0.4401|0.115|0.843|0.042|RT @HamiltonElector: RT The only thing that matters now is educating EVERYONE that Donald Trump is not President yet. He has not won. #Dec1
SAGEIntl66|edition|-0.4767|0.237|0.763|0.0|Closing ranks on Trump... dangerous times ahead for the US. https://t.co/aPbGIjerTY
AntonioCabeza_|TeenVogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
AntonioCabeza_|teenvogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
nofixedabode|jamestaranto|0.8124|0.0|0.72|0.28|"RT @jamestaranto: ""If facts become a point of debate, the very definition of freedom will be called into question."" Um, OK. https://t.co/12"
nofixedabode|t|0.8124|0.0|0.72|0.28|"RT @jamestaranto: ""If facts become a point of debate, the very definition of freedom will be called into question."" Um, OK. https://t.co/12"
MiaShaw|SenSanders|0.4767|0.08|0.691|0.229|"RT @SenSanders: I challenge Mr. Trump to tell the American people he'll keep his promises and veto cuts to Social Security, Medicare and Me"
MonicaFitz1|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
talene|tribelaw|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
talene|twitter|0.0|0.0|1.0|0.0|RT @tribelaw: Yup. That's exactly what he is. And now Trump tells us it's what he intends to be and do. https://t.co/6H5mmVEPkU
terrybrown5367|TeenVogue|0.0|0.0|1.0|0.0|Donald Trump Is Gaslighting America https://t.co/bKzYk9hIcU via @TeenVogue
terrybrown5367|linkis|0.0|0.0|1.0|0.0|Donald Trump Is Gaslighting America https://t.co/bKzYk9hIcU via @TeenVogue
C_BOYCE|quinncy|0.0|0.0|1.0|0.0|"RT @quinncy: I'm going to keep saying this. Trump needs his family around because he has Alzheimer's. They cover for him, keep him less anx"
sunlightwarden|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
sunlightwarden|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
daboogieman_|politico|0.0|0.0|1.0|0.0|"California elector files suit, joins anti-Trump Electoral College push https://t.co/a4L0WuDRM4 #hamiltonelectors #AuditTheVote #Resist"
honorverity|USA_Pragmatic1|0.3182|0.0|0.901|0.099|"RT @USA_Pragmatic1: @Khanoisseur @mms5048 That's 100% truth. Plus, the FACT Trump has been showing us for decades who he really is. https:/"
honorverity||0.3182|0.0|0.901|0.099|"RT @USA_Pragmatic1: @Khanoisseur @mms5048 That's 100% truth. Plus, the FACT Trump has been showing us for decades who he really is. https:/"
scoutinfinity|amjoyshow|-0.4404|0.132|0.868|0.0|"RT @amjoyshow: Scott Dworkin (@FUNDER) started #TrumpLeaks documenting hundreds of Trump's Russian ties, which the #FBI has denied or not r"
bluebonnetbunny|grumpyoldman418|0.5994|0.0|0.741|0.259|"RT @grumpyoldman418: Trump, Jr. Russians make up a pretty disproportionate cross-section of a lot of our assets,  https://t.co/ktNfyMSX9v"
bluebonnetbunny|linkis|0.5994|0.0|0.741|0.259|"RT @grumpyoldman418: Trump, Jr. Russians make up a pretty disproportionate cross-section of a lot of our assets,  https://t.co/ktNfyMSX9v"
Martina|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
Sailfish157|TomthunkitsMind|0.128|0.191|0.598|0.211|"RT @TomthunkitsMind: Trump supporters got played, will pay thru 401k's, foreclosures, predatory lending, higher gas prices, sale of public"
cocktailgurl17|Bluegirl_3|-0.7579|0.347|0.653|0.0|RT @Bluegirl_3: Teen Vogue editor pulls fire alarm on Trump gaslighting: He spun accusations of his falsehoods as bias https://t.co/czsi5
cocktailgurl17|t|-0.7579|0.347|0.653|0.0|RT @Bluegirl_3: Teen Vogue editor pulls fire alarm on Trump gaslighting: He spun accusations of his falsehoods as bias https://t.co/czsi5
Psalm11813|Jerusalem_Post|0.0|0.0|1.0|0.0|RT @Jerusalem_Post: Trump: Stay tuned for secretary of state https://t.co/n3HozAdVH9 #USElection https://t.co/mC8Sg8Japn
Psalm11813|jpost|0.0|0.0|1.0|0.0|RT @Jerusalem_Post: Trump: Stay tuned for secretary of state https://t.co/n3HozAdVH9 #USElection https://t.co/mC8Sg8Japn
seeker55|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: Trump: 'Nobody really knows' if #ClimateChange is real. Um... Apart from every scientist who works on the subject?! Idi
mmagoski01|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
parishatzi|forbes|0.0|0.0|1.0|0.0|Donald Trump's $100 Million Private Jet Features Gold-Plated (Nearly) Everything https://t.co/ppE3x8kiG2
Tweeting_Local|bloomberg|-0.34|0.179|0.821|0.0|business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/dYhaX42Jhk https://t.co/veYluNxQ2H
TroutlineCreek|VABVOX|0.0|0.0|1.0|0.0|"RT @VABVOX: 21) If #ElectoralCollege votes Trump regardless of the Putin/Russia connection, Congress can demand--must be in writing--a re-d"
throwinschade|Parker9_|0.875|0.0|0.643|0.357|RT @Parker9_: Funny how Trump supporters love to fly the flags of armies that got their asses kicked by Americans https://t.co/r4bN63AiuF
throwinschade|twitter|0.875|0.0|0.643|0.357|RT @Parker9_: Funny how Trump supporters love to fly the flags of armies that got their asses kicked by Americans https://t.co/r4bN63AiuF
eprophotog|funder|-0.2023|0.083|0.917|0.0|RT @funder: #TRUMPLEAKS:16 House Dems ask AG to investigate 25k bribe from Trump via Foundation for TrumpU#cnn #msnbc #AMJoy #cnnsotu #thi
mtighe15|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
bachic2|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
P1e2h7Patrick|twitter|-0.296|0.165|0.72|0.114|IRON: Trump vanguard of baby-boomers parents victory over fascism now introducing same 70 years after war WITH help https://t.co/Ll57tIIDxt
JodiMaxwell1|SenateGOP|-0.296|0.167|0.833|0.0|What RU hiding? @SenateGOP @HouseGOP @SpeakerRyan #RussiaHacking #russiahacker #russia #donthecon #trumplies https://t.co/HfZniSGvOX
JodiMaxwell1|bostonglobe|-0.296|0.167|0.833|0.0|What RU hiding? @SenateGOP @HouseGOP @SpeakerRyan #RussiaHacking #russiahacker #russia #donthecon #trumplies https://t.co/HfZniSGvOX
metroadlib|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
Beatromney|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: If Trump administration ends w/ Russia in control of Estonia and Latvia (directly or with his boys in charge), Putin's"
84Suburban|CNET|0.0|0.0|1.0|0.0|"RT @CNET: Larry Page, Tim Cook said to attend Donald Trump's tech summit https://t.co/6k7UqPrWJI https://t.co/1Bu6w6VOG3"
84Suburban|cnet|0.0|0.0|1.0|0.0|"RT @CNET: Larry Page, Tim Cook said to attend Donald Trump's tech summit https://t.co/6k7UqPrWJI https://t.co/1Bu6w6VOG3"
PaulieAbeles|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
PaulieAbeles|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
redge02|JoyAnnReid|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
redge02|twitter|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
djvrobin|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
djvrobin|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
arieella_|twitter|0.0|0.0|1.0|0.0|As if Trump isn't enough. As if 2016 hasn't been enough. https://t.co/J3TpBs28LX
xmssweetnessx|CathyLind2|0.0772|0.0|0.925|0.075|RT @CathyLind2: @transition2017 All I want for Christmas is to see @brunelldonald have a place in President Trump's administration.She's a
annwalker_13|SenSanders|0.2023|0.058|0.853|0.089|RT @SenSanders: Mr. Trump told working people he was on their side. Millions of us are going to demand that he keep his promise.
BlazeBerner|TrivWorks|0.0|0.0|1.0|0.0|"RT @TrivWorks: Trump: ""The Apprentice""Palin: ""Sarah Palin's Alaska""Rick Perry: ""Dancing with the Stars""This is the reality of our execu"
RussJensen5|FoxNews|0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
RussJensen5||0.0|0.0|1.0|0.0|"RT @FoxNews: .@JudgeJeanine: ""We have a new Pres.-elect. His name is Donald J. Trump. So move over, Barack. Move over, Hillary."" https://t."
TeaTraitors|Newyorker2212|-0.6808|0.286|0.714|0.0|@Newyorker2212 @DavidCornDC And Al Qaeda &amp; ISIS Deciding who attacks 1st since Trump ignoring Intel Reports.
melman456|SavageBiden|0.5719|0.0|0.709|0.291|@SavageBiden @miakhaIifa my reaction when Trump won the election... https://t.co/RTEmUJteOz
melman456|twitter|0.5719|0.0|0.709|0.291|@SavageBiden @miakhaIifa my reaction when Trump won the election... https://t.co/RTEmUJteOz
smokeyvera|SocialPowerOne1|0.0|0.0|1.0|0.0|"RT @SocialPowerOne1: The FBI Just Got Sued, And It Could Lead to Trumps Impeachment https://t.co/KASI7FtG93"
smokeyvera|occupydemocrats|0.0|0.0|1.0|0.0|"RT @SocialPowerOne1: The FBI Just Got Sued, And It Could Lead to Trumps Impeachment https://t.co/KASI7FtG93"
melindacasino|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
KirbAnne|20committee|0.2023|0.0|0.924|0.076|RT @20committee: Trump's refusal to admit that Russia was behind election games is forcing his cabinet nominees to lie publicly in ways the
bartelmoose|thehill|-0.6794|0.227|0.773|0.0|"@thehill ""Biden: Trump ran ""most vicious"" campaign I've ever seen"" ... Hillary's Campaign was equally as vicious, Joe ... @JoeBiden @VP"
BlueSpiderwort|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
BlueSpiderwort||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
joelderfner|annehelen|0.4767|0.063|0.791|0.146|RT @annehelen: Trump views his presidency as a narrative w/rising and falling action; note to journalists that he loves it when others do a
furngals2|NewtTrump|0.5267|0.0|0.861|0.139|"RT @NewtTrump: Newt explains Trump's MASTERFUL winning Twitter strategy ""If you don't give the media a rabbit to chase each day, they'll in"
pollomaldonado|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
pollomaldonado|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
bhendricks72013|twitter|0.0|0.0|1.0|0.0|"That, in and of itself, is enough reason to keep Trump out of the White House #hamiltonelectors https://t.co/KFueTJlthg"
JoelVanderWerf|DanRather|0.0|0.0|1.0|0.0|RT @DanRather: The question now is whether this will be a Trump Putin Administration or a Putin Trump Administration? https://t.co/PF20Xo89
JoelVanderWerf|t|0.0|0.0|1.0|0.0|RT @DanRather: The question now is whether this will be a Trump Putin Administration or a Putin Trump Administration? https://t.co/PF20Xo89
RobertA87413263|jmaboshie|0.8573|0.165|0.482|0.354|"RT @jmaboshie: Im Vladimir, i stole the election for #Trump but I let Hillary win the popular vote. I forgot to rig that part. My bad. Won'"
ToddDomke|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/U1KFDsn1Mf https://t.co/Z21lnE9BwB
ToddDomke|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/U1KFDsn1Mf https://t.co/Z21lnE9BwB
girishglg|kausmickey|0.4201|0.0|0.859|0.141|"RT @kausmickey: ""Nobody voted for [Trump] because they wanted him to be more like Bush on immigration."" https://t.co/BcShCvQBdg"
girishglg|conservativereview|0.4201|0.0|0.859|0.141|"RT @kausmickey: ""Nobody voted for [Trump] because they wanted him to be more like Bush on immigration."" https://t.co/BcShCvQBdg"
VorheesBev|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
mrapier|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
sanzimm|JuddLegum|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
sanzimm|medium|0.0|0.0|1.0|0.0|"RT @JuddLegum: 9. Anyway, this is who is advising Trump https://t.co/oRUPSkz7NV"
Brentm_5|TrumpNewMedia|-0.5147|0.237|0.64|0.123|RT @TrumpNewMedia: Having a #Traitor like @MittRomney as SOS would be a BETRAYAL! @realDonaldTrump @IvankaTrump @EricTrump @DonaldJTrumpJr
Rumky6|Will_Bunch|-0.7149|0.239|0.761|0.0|"RT @Will_Bunch: Worse than Watergate? Russia hacking is massive cloud over Trump presidency, and America. What caused this big mess? https:"
jackhenrynola|funder|-0.6808|0.248|0.752|0.0|"RT @funder: Breaking: We are filing complaints for treason tmrw on Trump, McConnell, Giuliani &amp; James Comey.#DworkinReport #TrumpLeaks Ru"
NickKilstein|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
cmalocksmith|nytimesworld|0.0|0.0|1.0|0.0|"RT @nytimesworld: What if ""North Korea offers to Donald Trump that there is a lot of real estate that he can develop in North Korea""? https"
Only4RM|EdSkipper|-0.6448|0.249|0.659|0.093|"RT @EdSkipper: Just as FYI - know SO MANY white middle class ""Christians"" still in rage and grief over Trump @Only4RM @missb62"
MarcLajambe|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Tea4gunsSC|twitter|-0.2057|0.232|0.768|0.0|We'll see I'm not a trump supporter https://t.co/z2Kp9BHTQy
lucas460|jrobertoacosta1|0.0|0.0|1.0|0.0|"RT @jrobertoacosta1: Por cuenta de incertidumbre por Trump, Mxico nos iguala en ""virreinato"" de Bonos mas riesgosos en mercados globales h"
oneinatree|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: US Senators letter to Senate leaders-investigate Trump for Russian espionage#cnn #msnbc #AMJoy #cnnsotu #thiswee
WilliamSnowHume|3NovicesChennai|-0.4019|0.197|0.803|0.0|"@3NovicesChennai Everyone should reject it, until the evidence is public. #CIA_Star_Chamber  https://t.co/ej1ykj3irM"
WilliamSnowHume|cnn|-0.4019|0.197|0.803|0.0|"@3NovicesChennai Everyone should reject it, until the evidence is public. #CIA_Star_Chamber  https://t.co/ej1ykj3irM"
kateb722|TrumpSuperPAC|-0.9106|0.435|0.565|0.0|RT @TrumpSuperPAC: Proof @CNN's #FakeNews. Watch stadium's reaction to hearing President-Elect TRUMP arrived! Racists? Nazis? Hell No!! htt
ndylan1|NormEisen|0.595|0.101|0.668|0.231|"RT @NormEisen: Wow, Trump has just 41% approval (vs 72 at this pt 4 Obama) with 65% concerned that his business ties CONFLICT. https://t.co"
ndylan1|t|0.595|0.101|0.668|0.231|"RT @NormEisen: Wow, Trump has just 41% approval (vs 72 at this pt 4 Obama) with 65% concerned that his business ties CONFLICT. https://t.co"
BRTTVNY_|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
VijayKulkarnii|Forbes|0.0|0.0|1.0|0.0|RT @Forbes: Take a look inside Trump's $100 million private jet: https://t.co/CfrvKeExGp https://t.co/Ar3DfhnLOH
VijayKulkarnii|forbes|0.0|0.0|1.0|0.0|RT @Forbes: Take a look inside Trump's $100 million private jet: https://t.co/CfrvKeExGp https://t.co/Ar3DfhnLOH
BarusArus|FortuneMagazine|0.4215|0.0|0.843|0.157|RT @FortuneMagazine: Netanyahu says he hopes to work with Trump to undo Iran deal https://t.co/NXEDvuTJQC https://t.co/xeuV1vVKtu
BarusArus|fortune|0.4215|0.0|0.843|0.157|RT @FortuneMagazine: Netanyahu says he hopes to work with Trump to undo Iran deal https://t.co/NXEDvuTJQC https://t.co/xeuV1vVKtu
Pink22Karen|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
Pink22Karen|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
mama2fluffs|kylegriffin1|-0.6124|0.2|0.8|0.0|RT @kylegriffin1: Two longtime ethics experts argue Trump's biz conflicts are so big it should affect how the Electoral College votes: http
hsjr33|WayneDupreeShow|-0.4767|0.171|0.829|0.0|RT @WayneDupreeShow: Rep. Tulsi Gabbard Says Democrats Wrong To Bash Trump For Retired General Picks https://t.co/62oDMIBBmO
hsjr33|newsninja2012|-0.4767|0.171|0.829|0.0|RT @WayneDupreeShow: Rep. Tulsi Gabbard Says Democrats Wrong To Bash Trump For Retired General Picks https://t.co/62oDMIBBmO
KarenOggs|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
KarenOggs|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
ausyj|riotbookshelf|-0.7351|0.289|0.647|0.065|RT @riotbookshelf: I outraged my relatives by 'generalising' Trump voters. Fact remains they all voted for a white supremacist perpetrator
MrsRothenberg|TheDemocrats|0.5514|0.0|0.818|0.182|RT @TheDemocrats: Are you:- A woman?- Under 26?Do you:- Have a pre-existing condition?- Live?- Breathe?Obamacare helps you. Don't le
remmkm|JohnRMoffitt|-0.2023|0.116|0.8|0.084|"RT @JohnRMoffitt: Well, as #Trump famously said, ""What's the point of having all these nuclear weapons if we don't use them?"" https://t.co/"
remmkm|t|-0.2023|0.116|0.8|0.084|"RT @JohnRMoffitt: Well, as #Trump famously said, ""What's the point of having all these nuclear weapons if we don't use them?"" https://t.co/"
Tull007|JuddLegum|0.128|0.0|0.897|0.103|RT @JuddLegum: 2. He's also a leading contender to be Deputy Secretary of State https://t.co/oRUPSkz7NV
Tull007|medium|0.128|0.0|0.897|0.103|RT @JuddLegum: 2. He's also a leading contender to be Deputy Secretary of State https://t.co/oRUPSkz7NV
anastasialie83|twitter|-0.3291|0.11|0.89|0.0|"If it's secret, how do u know?Also, you're behind. It's an attempt 2 keep trump out of office. I hate him, but I https://t.co/UyHDdEWfb9"
eduardoinalbion|Evan_McMullin|-0.1027|0.129|0.759|0.112|"RT @Evan_McMullin: Trump encouraged Russian subversion of our democracy then denied its occurrence despite CIA evidence, while preparing to"
BrunoG_Gallo|borjaechevarria|0.0|0.0|1.0|0.0|RT @borjaechevarria: A private club in Palm Beach is the Trump company that requested the most U.S. work visas for foreign nationals https:
mapnotes|dailynewsbin|0.0|0.0|1.0|0.0|https://t.co/EPXOv9ogq7
NettaBear13|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
julie2too|nattie8859|0.0|0.0|1.0|0.0|"@nattie8859 @Vzladream @FoxNews That would be you and Trump, right. Keep your religion and I'll keep mine."
sanzimm|JuddLegum|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
sanzimm|medium|-0.3182|0.187|0.813|0.0|RT @JuddLegum: 8. Even the Fox News people were shocked https://t.co/oRUPSkz7NV
hknyemi|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Jillsey11|noamscheiber|-0.4215|0.141|0.859|0.0|RT @noamscheiber: Your next labor secretary insists Obamacare has caused a restaurant recession. The data insists the opposite https://t.co
Jillsey11|t|-0.4215|0.141|0.859|0.0|RT @noamscheiber: Your next labor secretary insists Obamacare has caused a restaurant recession. The data insists the opposite https://t.co
randomirish|theguardian|-0.0258|0.196|0.613|0.19|Intelligence figures fear Trump reprisals over assessment of Russia election role https://t.co/72QiRkZVjq
lspesq53_lsp|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
TovarRasputin|realDonaldTrump|0.4767|0.0|0.807|0.193|The words Trump &amp; Intelligence are orthogonal. (look that up @realDonaldTrump &amp; #trumpchumps) https://t.co/dNl6ietCn8
TovarRasputin|twitter|0.4767|0.0|0.807|0.193|The words Trump &amp; Intelligence are orthogonal. (look that up @realDonaldTrump &amp; #trumpchumps) https://t.co/dNl6ietCn8
iyamiyam|JohnFugelsang|-0.2263|0.087|0.913|0.0|RT @JohnFugelsang: Trump blocks #millionwomanmarch from Lincoln Memorial despite the fact that the LM is actually owned by Americans who pa
BusMinCommunity|bloomberg|-0.34|0.179|0.821|0.0|business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/T1cf5qQ0ZS https://t.co/RZrywZS6k2
8thhousegoddess|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
mattydubswack|StefanMolyneux|-0.5423|0.289|0.597|0.114|RT @StefanMolyneux: The Truth About Fake NewsRussia Hacked U.S. Election For Donald Trump? https://t.co/L1g8OJzXRr https://t.co/Oiww50IJSY
mattydubswack|youtube|-0.5423|0.289|0.597|0.114|RT @StefanMolyneux: The Truth About Fake NewsRussia Hacked U.S. Election For Donald Trump? https://t.co/L1g8OJzXRr https://t.co/Oiww50IJSY
AmericasImpetus|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
luvauntyruth|KellyAuCoin77|0.0|0.0|1.0|0.0|RT @KellyAuCoin77: Trump Picks El Chapo to Run D.E.A. https://t.co/U1kSzcRlA1 via @BorowitzReport
luvauntyruth|newyorker|0.0|0.0|1.0|0.0|RT @KellyAuCoin77: Trump Picks El Chapo to Run D.E.A. https://t.co/U1kSzcRlA1 via @BorowitzReport
tai_barron|_jackkrecidlo|0.4144|0.0|0.765|0.235|RT @_jackkrecidlo: This snow is so white it supports trump
margab18|HuffPostPol|0.0|0.0|1.0|0.0|"Donald Trump says it is ""ridiculous"" to say Russia intervened in the election on his behalf. https://t.co/OMmJXNzNIC via @HuffPostPol"
margab18|huffingtonpost|0.0|0.0|1.0|0.0|"Donald Trump says it is ""ridiculous"" to say Russia intervened in the election on his behalf. https://t.co/OMmJXNzNIC via @HuffPostPol"
thebobbyb|politicususa|0.3182|0.105|0.718|0.177|Hell-Surrogate = KushnerTrump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests via @politicususa https://t.co/BjrZayhcT6
thebobbyb|politicususa|0.3182|0.105|0.718|0.177|Hell-Surrogate = KushnerTrump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests via @politicususa https://t.co/BjrZayhcT6
tray24u1|bfraser747|0.0|0.0|1.0|0.0|"RT @bfraser747: ""We have a new PresElect. His name is Donald J. Trump. So move over, Barack Move over Hillary"" AMEN @JudgeJeaninehttps:/"
apwriter|twitter|0.5562|0.0|0.841|0.159|Have fun at the pump Trumpkins! Mr. Exxon means oil futures up 5% tonight already. U was robbed. #russia #trump https://t.co/JDWaFNTTWn
PHLBizDPoncet|kurteichenwald|0.5574|0.0|0.847|0.153|"RT @kurteichenwald: If Trump started getting praise 4  appointments from ISIS, do you think Fox News would start running stories about how"
michaelpsycho|YourAnonCentral|-0.4939|0.144|0.856|0.0|"RT @YourAnonCentral: Steal this: Open Call for mobilization against the inauguration of Donald #Trump on January 20, 2017 #DisruptJ20  http"
clotfelter11|MichaelGaree|-0.5267|0.204|0.739|0.057|"RT @MichaelGaree: Something comrade Trump's inner circle might want to consider: If he's charged with treason, guess who becomes co-conspir"
BusMinCommunity|twitter|0.6249|0.062|0.705|0.232|business: RT bpolitics: Trump says his support for the One-China policy will hinge on cutting a better deal on tra https://t.co/fr5StJfUfp
DebbieW36246900|JuddLegum|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
DebbieW36246900|t|0.4588|0.0|0.87|0.13|"RT @JuddLegum: 4. Bolton called it a ""false flag,"" which is a favorite term of InfoWars, the people who brought you pizzagate https://t.co/"
BiasedGirl|twitter|0.0|0.0|1.0|0.0|You know President-elect Trump is going to be tweeting about this... https://t.co/ZKymGISMXs
VlDEOSTARK|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
maruhkati|pixelatedboat|-0.4585|0.167|0.833|0.0|RT @pixelatedboat: I read the 12th Amendment and technically neither Clinton nor Trump won the election: https://t.co/fKieKK3fEH
maruhkati|twitter|-0.4585|0.167|0.833|0.0|RT @pixelatedboat: I read the 12th Amendment and technically neither Clinton nor Trump won the election: https://t.co/fKieKK3fEH
PatVPeters|DailyCaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
PatVPeters|dailycaller|0.34|0.0|0.862|0.138|RT @DailyCaller: Sen. Tim Scott Lays Out Plan For Trump To Engage Black Communities https://t.co/uXRD9iaGsd https://t.co/dOJr3MhDaF
lyz_estrada|GOPjenna|-0.5859|0.219|0.704|0.078|RT @GOPjenna: It's obvious u guys r upset cuz your attempt w the Reince/Romney deal failed. Trump &amp; his army of loyalists will ALWAYS outsm
didi8367|johnpavlovitz|-0.0725|0.055|0.945|0.0|RT @johnpavlovitz: I wouldn't have to talk so much about Donald Trump if you didn't say so little. I won't apologize for being fully oppose
Froghorn2016|Lrihendry|0.1275|0.113|0.756|0.13|RT @Lrihendry: While shopping 2day I overheard a conv with group saying isn't it great we can say Merry Christmas again &amp; not be afraid! WO
Carlapaul18|V_of_Europe|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
Carlapaul18|thegatewaypundit|-0.0772|0.253|0.553|0.194|RT @V_of_Europe: Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
chimeraelf|JordanChariton|-0.4404|0.162|0.838|0.0|"RT @JordanChariton: This is BEYOND THE PALE, even for @realDonaldTrump. Dems need to block this https://t.co/LnniEBcwnu"
chimeraelf|nbcnews|-0.4404|0.162|0.838|0.0|"RT @JordanChariton: This is BEYOND THE PALE, even for @realDonaldTrump. Dems need to block this https://t.co/LnniEBcwnu"
WizardOfOsrin|DenbrotS|0.0|0.0|1.0|0.0|RT @DenbrotS: @NancyPelosi @blueskymountain @HouseGOP Of course Trump will stiff the miners. He's silent.
ThelmaOAgyekum|CNN|-0.4215|0.135|0.865|0.0|"RT @CNN: This county voted Democrat for 144 years. But in 2016, Donald Trump broke that streak https://t.co/cFNxi10sCK https://t.co/dhxrTti"
ThelmaOAgyekum|cnn|-0.4215|0.135|0.865|0.0|"RT @CNN: This county voted Democrat for 144 years. But in 2016, Donald Trump broke that streak https://t.co/cFNxi10sCK https://t.co/dhxrTti"
WkndGirl|TeaPainUSA|0.0516|0.086|0.822|0.092|RT @TeaPainUSA: Is there any doubt left as to why Donald Trump won't release his tax returns?  Red Don needs to come clean or concede.  #Tr
THEJEDEYE1|latimes|-0.4019|0.172|0.828|0.0|RT @latimes: The obscure constitutional provision that could be trouble for Trump https://t.co/yv5pTs6c32 https://t.co/4ZLRELxfbs
THEJEDEYE1|latimes|-0.4019|0.172|0.828|0.0|RT @latimes: The obscure constitutional provision that could be trouble for Trump https://t.co/yv5pTs6c32 https://t.co/4ZLRELxfbs
abbeysbooks|JSavoly|-0.4019|0.137|0.863|0.0|RT @JSavoly: Trump Gives The Electoral College Reason To Reject Him During Fox News Interview #StollenElection #ComradeTrump  https://t.co/
abbeysbooks|t|-0.4019|0.137|0.863|0.0|RT @JSavoly: Trump Gives The Electoral College Reason To Reject Him During Fox News Interview #StollenElection #ComradeTrump  https://t.co/
cnewionlpn|saladinahmed|-0.6704|0.29|0.71|0.0|RT @saladinahmed: TRUMP'S CABINET is an anagram of 'TIS BUT CRAP MEN
PatPatojson|Corporatocrazy|-0.5594|0.18|0.82|0.0|"RT @Corporatocrazy: So the CIA leaks fake news to media and then wonders why Trump doesn't want to attend daily ""intelligence"" briefing! SM"
ShonaLovesTrump|snip|0.7269|0.0|0.596|0.404|LETTER TO THE EDITOR: Obama responsible for Donald Trump win https://t.co/xWjVHEEn1D
c4trends|twitter|0.0|0.0|1.0|0.0|"what does #Bill Gates, #Ma and John #Doerr know that #Trump doesn't? https://t.co/EpFv1z9lus"
SusanCarver19|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
greenwonk|transportgooru|0.25|0.0|0.882|0.118|The golden age of US #infrastructure - will Trump's vision come even close? @transportgooru @CoryBooker @SenSanders https://t.co/4K0FFlERDK
greenwonk|twitter|0.25|0.0|0.882|0.118|The golden age of US #infrastructure - will Trump's vision come even close? @transportgooru @CoryBooker @SenSanders https://t.co/4K0FFlERDK
mattbaumanNYC|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
pettywap7teen38|MichaelSkolnik|-0.4588|0.125|0.875|0.0|RT @MichaelSkolnik: Many Republicans are going to have a rude awakening when they finally realize what we all have known. Trump is putting
harley_gernand|mikandynothem|0.5859|0.0|0.826|0.174|"RT @mikandynothem: President-elect Donald Trump defied all odds to win Presidency. We are looking at next Reagan, America. Perhaps...even g"
HoosierMum|Will_Bunch|-0.7149|0.239|0.761|0.0|"RT @Will_Bunch: Worse than Watergate? Russia hacking is massive cloud over Trump presidency, and America. What caused this big mess? https:"
websterwakeemup|Lee_in_Iowa|-0.1531|0.191|0.674|0.135|"@Lee_in_Iowa @adirado29 If lies and innuendo can win an election for Trump, who has lied repeatedly,the nation turns it's head in disbelief."
theshoewife|NBCNews|0.0516|0.145|0.661|0.194|RT @NBCNews: A slap in the face. That's how intelligence agencies see Trump's rejection of findings on Russia https://t.co/k6QZxwjtem https
theshoewife|nbcnews|0.0516|0.145|0.661|0.194|RT @NBCNews: A slap in the face. That's how intelligence agencies see Trump's rejection of findings on Russia https://t.co/k6QZxwjtem https
ShonaLovesTrump|snip|0.0|0.0|1.0|0.0|Donald Trump should meet with King Hamad of Bahrain https://t.co/gYvaaoY5Fp
sadhana456|kylegriffin1|-0.5267|0.145|0.855|0.0|"RT @kylegriffin1: Watergate reporter Carl Bernstein: 'Nixon was nothing, in terms of lying, compared to what we've seen from Trump.' https:"
venead12|ecotalvora|0.0|0.0|1.0|0.0|RT @ecotalvora: Segn DEA Farc @FARC_EPueblo es eslabn d  narcotrfico pese  negociaciones d paz #InformeOtlvora #Colombia https://t.co
venead12|t|0.0|0.0|1.0|0.0|RT @ecotalvora: Segn DEA Farc @FARC_EPueblo es eslabn d  narcotrfico pese  negociaciones d paz #InformeOtlvora #Colombia https://t.co
hgreenberg1|TeaPainUSA|0.6808|0.0|0.772|0.228|RT @TeaPainUSA: Trump's tryin' to save America.  The fewer security briefings he receives the fewer he has to forward to Putin.https://t.
theonlyadult|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
TroncaleJoseph|_News_Trump|-0.4336|0.265|0.617|0.118|@_News_Trump #AbandonHopeAllYeWhoEnterSafeSpaces. You are sheep inviting slaughter. You are so unsafe. The irony is pathetic.
lanatwotwo|politicususa|0.3182|0.09|0.758|0.152|RT @politicususa: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests via @politicususa https://t.co/IKDOxKghqQ #p2 #c
lanatwotwo|politicususa|0.3182|0.09|0.758|0.152|RT @politicususa: Trump Surrogate Calls on FBIs Comey to Crackdown on Peaceful Protests via @politicususa https://t.co/IKDOxKghqQ #p2 #c
brloggins3412|eddiespike|-0.7003|0.236|0.764|0.0|"RT @eddiespike: Dont give a damn if your Dem or Rep, Trump or Clinton, just stop whining. Work toward positve change or just quit your endl"
Emmita17E|DrEstella|0.0|0.0|1.0|0.0|"RT @DrEstella: Senator #HarryRead asks CIA to lie to @realDonaldTrump ""Give Trump ""Fake"" INTEL BRIEFINGS!""  #SundayMorning #WeareTrump #Tru"
VeroPArtist|ABFalecbaldwin|0.9057|0.13|0.307|0.563|Awesome! @ABFalecbaldwin won best guest actor for #SNL playing stupid #trump !!  #CriticsChoiceAwards
Pellagios|_Makada_|-0.296|0.115|0.826|0.06|"RT @_Makada_: President-Elect Trump: It's ridiculous to say Russia intervened in the election, I think it's just another excuse. We had a m"
maegabby49|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
maegabby49|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
kldreams61|NewtTrump|0.5267|0.0|0.861|0.139|"RT @NewtTrump: Newt explains Trump's MASTERFUL winning Twitter strategy ""If you don't give the media a rabbit to chase each day, they'll in"
BruinsRocknRule|hectormorenco|-0.6369|0.284|0.608|0.108|RT @hectormorenco: Trump should repeal and replace Obama Care for no other reason than to trash arrogant &amp; obnoxious Obama's signature dome
AnnH1958|dailycaller|0.0|0.0|1.0|0.0|https://t.co/Tfh8PwLgrL
MarkStemen|theonlyadult|0.6249|0.0|0.812|0.188|"RT @theonlyadult: If you didn't vote for Hillary, you voted for Trump. The rest is just garbage words salad to feel better about helping a"
ReclaimDawgs|mitchellvii|-0.5994|0.214|0.786|0.0|RT @mitchellvii: When is the Media going to learn that Americans no longer give a damn what they say about Trump?
carolefeuerman|StoneSculptorJN|0.0|0.0|1.0|0.0|RT @StoneSculptorJN: Donald Trump Wants To Abolish The Federal Reserve  https://t.co/Bs3w4RAXCZ
carolefeuerman|whydontyoutrythis|0.0|0.0|1.0|0.0|RT @StoneSculptorJN: Donald Trump Wants To Abolish The Federal Reserve  https://t.co/Bs3w4RAXCZ
dogmotto|Joyce_Karam|-0.8176|0.309|0.691|0.0|RT @Joyce_Karam: There's an attack on Church in Egypt;Terror in Istanbul; ISIS took Palmyra; CIA alarm on Russia.But #Trump is attacking NB
instinctnaturel|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
waltercwawalter|halconada|0.0|0.0|1.0|0.0|RT @halconada: La noticia del da: el gobierno de EEUU afirma que hackers de Rusia ayudaron  a Trump durante la campaa electoral: https://
waltercwawalter||0.0|0.0|1.0|0.0|RT @halconada: La noticia del da: el gobierno de EEUU afirma que hackers de Rusia ayudaron  a Trump durante la campaa electoral: https://
Aubrey_Gayle|gollum1419_g|0.0516|0.145|0.7|0.155|"RT @gollum1419_g: As Trump again attacks CIA, former intelligence officers expect retaliation https://t.co/RmPY9nxbFP #Trump #Corruption #W"
Aubrey_Gayle|dailykos|0.0516|0.145|0.7|0.155|"RT @gollum1419_g: As Trump again attacks CIA, former intelligence officers expect retaliation https://t.co/RmPY9nxbFP #Trump #Corruption #W"
Barkforlove1|twitter|-0.3382|0.194|0.684|0.121|So that means Bolton is a sure thing for team trump. Conspiracy theory nutters unite! https://t.co/t6cf8gY3j6
msjbe20a|NPR|0.0|0.0|1.0|0.0|Via @NPR: CIA Concludes Russian Interference Aimed To Elect Trump https://t.co/d8HD0puSHX
msjbe20a|npr|0.0|0.0|1.0|0.0|Via @NPR: CIA Concludes Russian Interference Aimed To Elect Trump https://t.co/d8HD0puSHX
realdadinstands|joanwalsh|0.0|0.0|1.0|0.0|@joanwalsh @HistoryInPics trump is going to do this right?  #fakenews
wotshaking|whatshaking|0.0|0.0|1.0|0.0|Trump: Nobody really knows if climate change isreal https://t.co/wyeHm7BWnX
gavoweb|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Tull007|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
Tull007|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
1549321s|liberalsociety|0.0|0.0|1.0|0.0|"Liz Warren Just Made Epic Federal Move Against Trumps Corruption, Holy Sh*t [Details] - https://t.co/mh8EAKk8Vp"
SashaMichael22|youtube|0.4019|0.0|0.769|0.231|https://t.co/a7pcf5v3B8#BREAKING #trump #BernieSanders #share #RogueOne #Strictly Trump benefitted from Sanders.
Psalm11813|Jerusalem_Post|0.0|0.0|1.0|0.0|RT @Jerusalem_Post: Trump says US not necessarily bound by 'one China' policy https://t.co/3NoDj12Qjw #BreakingNews
Psalm11813|jpost|0.0|0.0|1.0|0.0|RT @Jerusalem_Post: Trump says US not necessarily bound by 'one China' policy https://t.co/3NoDj12Qjw #BreakingNews
MikeHighley1|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
ConHaterFromAB|Gizmodo|-0.4939|0.314|0.686|0.0|@Gizmodo Trump should be jailed. Lock him up
2ndsights|WillBlackWriter|0.3182|0.0|0.897|0.103|RT @WillBlackWriter: Please tweet and ask your followers to tweet this Vine of Donald Trump asking Russia to hack Clinton. #Treasonhttps
JkFlower60|pierre|0.1027|0.104|0.741|0.156|"RT @pierre: Before Trump: ""You're entitled to your opinion, but you're not entitled to your own facts."" Now: there are no facts. https://t."
JkFlower60||0.1027|0.104|0.741|0.156|"RT @pierre: Before Trump: ""You're entitled to your opinion, but you're not entitled to your own facts."" Now: there are no facts. https://t."
Donna_DHKBB|SheWhoVotes|0.7297|0.0|0.679|0.321|RT @SheWhoVotes: HUGE: Paul Manafort's mini-me in Ukraine is a (former?) Russian intelligence operative: https://t.co/1cNnfu3jGX #TrumpPuti
Donna_DHKBB|politico|0.7297|0.0|0.679|0.321|RT @SheWhoVotes: HUGE: Paul Manafort's mini-me in Ukraine is a (former?) Russian intelligence operative: https://t.co/1cNnfu3jGX #TrumpPuti
magresta|twitter|0.5267|0.0|0.726|0.274|"And Trump, Bannon et al full of passionate intensity. https://t.co/sFexKXwQdx"
AnitaStubbs|activist360|0.0|0.0|1.0|0.0|RT @activist360: REPORT: Obsequious a**-kisser Trump's had his head up the colorectal cavities of Russian oligarchs for three decades https
ProAssad|DPRK_News|0.7184|0.0|0.739|0.261|"RT @DPRK_News: Donald Trump foreign minister Rex Tillerson receives Russian Federation Medal of Friendship, reserved for obedient slaves of"
melodyhultgren|billyeichner|0.6486|0.125|0.554|0.321|"RT @billyeichner: Democrats deserve better than Trump. Republicans deserve better than Trump. All Americans deserve better than this lying,"
RepublicanRehab|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
Hitokiri1|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
Hitokiri1|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
AyeAtheist|CBSNews|0.0|0.0|1.0|0.0|"RT @CBSNews: After seeing some of it curtailed post-Ferguson, police expect Trump to step up surplus military gear availability https://t.c"
AyeAtheist||0.0|0.0|1.0|0.0|"RT @CBSNews: After seeing some of it curtailed post-Ferguson, police expect Trump to step up surplus military gear availability https://t.c"
rachmanworks|paddyhirsch|0.6597|0.0|0.748|0.252|"RT @paddyhirsch: Trump waves carrot and stick at US firms ""Number one were going to treat them well, and number two there are going to be"
freedfried|mikandynothem|0.3802|0.088|0.767|0.146|RT @mikandynothem: Ruth Bader Ginsburg said she would resign if Trump won. Hit the road lady! That will give Trump even more Conservatives
hawaiianlove68|JSavoly|0.0|0.0|1.0|0.0|RT @JSavoly: Chris Christie Reportedly Told Trump To Take His Cabinet Positions And Shove Em #StollenElection #ComradeTrump  https://t.co/
hawaiianlove68|t|0.0|0.0|1.0|0.0|RT @JSavoly: Chris Christie Reportedly Told Trump To Take His Cabinet Positions And Shove Em #StollenElection #ComradeTrump  https://t.co/
ramix365|cnn|-0.2023|0.265|0.735|0.0|Donald Trump's controversial 'Apprentice' role https://t.co/z0TW0iUFdk
yanachoen|jasoninthehouse|0.0|0.0|1.0|0.0|.@jasoninthehouse: Investigate Trump's finances https://t.co/Su23AI0e9Z @moveon
yanachoen|petitions|0.0|0.0|1.0|0.0|.@jasoninthehouse: Investigate Trump's finances https://t.co/Su23AI0e9Z @moveon
mollylmaguire|azmoderate|-0.1779|0.261|0.541|0.198|RT @azmoderate: Did Donald Trump Commit Treason? https://t.co/66dDzAbKnS
mollylmaguire|nbcnews|-0.1779|0.261|0.541|0.198|RT @azmoderate: Did Donald Trump Commit Treason? https://t.co/66dDzAbKnS
petrified_syrup|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
TheJonFerns|MockDraftHQ|0.4404|0.0|0.805|0.195|RT @MockDraftHQ: #Trump Supporters Vandalize NFL Player's Home With Slurs #MAGA https://t.co/nBWudDFzJV #donaldtrump
TheJonFerns|mockdrafthq|0.4404|0.0|0.805|0.195|RT @MockDraftHQ: #Trump Supporters Vandalize NFL Player's Home With Slurs #MAGA https://t.co/nBWudDFzJV #donaldtrump
IndiaJenkins1|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
bdanaher17|linkis|0.2732|0.0|0.811|0.189|Rick Perry a leading candidate for U.S. energy post: source https://t.co/Xwhwq1IZ9k
RoughAcres|lauriecrosswell|0.0|0.0|1.0|0.0|RT @lauriecrosswell: Paul Ryan's transformation into a TrumpPence Stepford husband took less time than Trump's tax audit. #60Minutes
lapierre_george|linkis|0.2577|0.0|0.873|0.127|GOP SENATORS CHALLENGE #Trump on secretary of state prospect's Russia ties - FOX NEWS https://t.co/D9F4zRH9YT Hotpage_News
ravenhairgirl|helenmaryme|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
ravenhairgirl|twitter|0.0|0.0|1.0|0.0|RT @helenmaryme: #BadNewsFromTheInternet Trump still hasn't deleted his Twitter account https://t.co/j6Y1MpOb4x
ajordan1911|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
ajordan1911|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
SKCfan1|EnviroNews|0.4215|0.098|0.684|0.218|RT @EnviroNews: #Trump Portfolio Riddled w/ Oil Stocks - Conflict of Interest for Him to Sign Energy Bills? https://t.co/jKKyuJOZaT https:/
SKCfan1|environews|0.4215|0.098|0.684|0.218|RT @EnviroNews: #Trump Portfolio Riddled w/ Oil Stocks - Conflict of Interest for Him to Sign Energy Bills? https://t.co/jKKyuJOZaT https:/
NateInPhilly|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
tarpsy|FeministaJones|-0.5106|0.18|0.82|0.0|RT @FeministaJones: Hey. I'm gonna be on c-span tomorrow morning talking about poverty in a Trump administration
PennyLDuncan|starknightz|0.0|0.0|1.0|0.0|"RT @starknightz: U.S Intel community is stumped: ""What to do with a Trump who doesn't buy our BS?"" https://t.co/84HTKFw7NN #TrumpTrain #Pre"
PennyLDuncan|sott|0.0|0.0|1.0|0.0|"RT @starknightz: U.S Intel community is stumped: ""What to do with a Trump who doesn't buy our BS?"" https://t.co/84HTKFw7NN #TrumpTrain #Pre"
juanrentsnow88|Judgenap|0.925|0.0|0.309|0.691|@Judgenap GOD BLESS AMERICAGOD BLESS DONALD TRUMPGOD BLESS.  NAPOLITANOMERRY CHRISTMAS
mercedesfduran|nick_dacosta|0.5859|0.0|0.648|0.352|RT @nick_dacosta: Brilliant Norwegian cartoon on #Trump https://t.co/H4amqJQCFe
mercedesfduran|twitter|0.5859|0.0|0.648|0.352|RT @nick_dacosta: Brilliant Norwegian cartoon on #Trump https://t.co/H4amqJQCFe
MikeAndy128|starfirst|0.7351|0.0|0.721|0.279|"RT @starfirst: President Obamas approval rating hits new high, Donald Trumps approval rating in toilet https://t.co/sejTKFqwav via @daily"
MikeAndy128|dailynewsbin|0.7351|0.0|0.721|0.279|"RT @starfirst: President Obamas approval rating hits new high, Donald Trumps approval rating in toilet https://t.co/sejTKFqwav via @daily"
Witchy_99|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
DcLincoln761|activist360|-0.8316|0.291|0.709|0.0|"RT @activist360: THIS IS TODAY'S GOP: Trump has normalized racism, hate, bigotry and misogyny  and now Mitch McConnell is normalizing trea"
ChrisCassara|JINCHURIKl|-0.0772|0.075|0.925|0.0|RT @JINCHURIKl: when trump says hes gonna build a wall but you have a trick up your sleeve https://t.co/tdvu1qPqUM
ChrisCassara|vine|-0.0772|0.075|0.925|0.0|RT @JINCHURIKl: when trump says hes gonna build a wall but you have a trick up your sleeve https://t.co/tdvu1qPqUM
rjpierce|RobertKennedyJr|0.0|0.0|1.0|0.0|RT @RobertKennedyJr: The #USDeptofEnergy expects wind to generate 10% of Americas electricity by 2020 https://t.co/CxdsISINzO
rjpierce|fortune|0.0|0.0|1.0|0.0|RT @RobertKennedyJr: The #USDeptofEnergy expects wind to generate 10% of Americas electricity by 2020 https://t.co/CxdsISINzO
kramkardam|K_J_Marks|0.4404|0.129|0.597|0.274|"@K_J_Marks they're like Trump supporters. If they kiss the tram's ass hard enough they'll like them back, but deep inside they know..."
Holleewood92|TeenVogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
Holleewood92|teenvogue|0.4019|0.11|0.705|0.185|RT @TeenVogue: Donald Trump is gas lighting America and deliberately undermining the very foundation of our freedom https://t.co/M00m2yjuly
djvrobin|asamjulian|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
djvrobin|twitter|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
lapierre_george|linkis|0.0|0.0|1.0|0.0|#TRUMP LASHES OUT at NBC News on Twitter - THE HILL https://t.co/W5VQGlvlwI Hotpage_News
ClassicShadoww|RuthHHopkins|0.5859|0.0|0.847|0.153|RT @RuthHHopkins: Russia helped Trump win. The CIA has confirmed this. The election is invalid. There's opinions &amp; there's facts. This is f
PrissiKrissi3|twitter|0.0|0.0|1.0|0.0|"I guess Trump, trumped them https://t.co/thCHkB2U65"
rojophotography|EW|0.0|0.0|1.0|0.0|Bryan Cranston Brings Back Walter White for 'SNL' Trump Sketch https://t.co/iwba2p69eG via @EW
rojophotography|ew|0.0|0.0|1.0|0.0|Bryan Cranston Brings Back Walter White for 'SNL' Trump Sketch https://t.co/iwba2p69eG via @EW
AZULCAMPEON10|JonRiley7|-0.4019|0.163|0.837|0.0|"RT @JonRiley7: Stop blaming those who took Trump ""literally but not seriously."" Don't tell me we shouldn't take candidates' policy proposal"
washburnt|JohnDelury|-0.7469|0.189|0.811|0.0|"RT @JohnDelury: Not to be alarmist, but when I asked what Beijing will do if Trump persists w Two China Policy, the answer was war https://"
washburnt||-0.7469|0.189|0.811|0.0|"RT @JohnDelury: Not to be alarmist, but when I asked what Beijing will do if Trump persists w Two China Policy, the answer was war https://"
namastaebitches|KellyannePolls|-0.1779|0.082|0.918|0.0|@KellyannePolls @Newsweek anyone who slept with both Fred Thompson AND Donald Trump can NOT be taken seriously #homewrecker. #whore #badmom
SteveGarard|2ALAW|0.4048|0.0|0.786|0.214|RT @2ALAW: Isn't Christmas A Little More Special This Year? #MAGA#Trump https://t.co/o4QjFjrFEi
SteveGarard|twitter|0.4048|0.0|0.786|0.214|RT @2ALAW: Isn't Christmas A Little More Special This Year? #MAGA#Trump https://t.co/o4QjFjrFEi
WkndGirl|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
WkndGirl||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
pas5974|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
Humanitarian66|twitter|0.0|0.0|1.0|0.0|Q: what does Trump the Fowl say?A: cuck cuck #MAGA https://t.co/8043V9NsLF
PoppeDoctor|FoxNews|-0.296|0.145|0.855|0.0|"RT @FoxNews: .@ericbolling: Trump to Stop 'Banksters', CEOs From 'Fooling' Average Americans https://t.co/MvCy3Ou08b https://t.co/Mq5RkPThrV"
PoppeDoctor|insider|-0.296|0.145|0.855|0.0|"RT @FoxNews: .@ericbolling: Trump to Stop 'Banksters', CEOs From 'Fooling' Average Americans https://t.co/MvCy3Ou08b https://t.co/Mq5RkPThrV"
Bnkr_Chk2|Seanbabydotcom|-0.743|0.294|0.615|0.091|RT @Seanbabydotcom: The BOP says 8.5% of prisoners are sex offenders. That fucking means a woman is 2.2 times safer in a federal prison tha
KimbyHuffy|amjoyshow|-0.3612|0.217|0.783|0.0|RT @amjoyshow: Blueprint for fighting Donald Trump https://t.co/GLMez1CsDU via @amjoyshow
KimbyHuffy|msnbc|-0.3612|0.217|0.783|0.0|RT @amjoyshow: Blueprint for fighting Donald Trump https://t.co/GLMez1CsDU via @amjoyshow
KittenMcKay|ericgarland|0.5719|0.0|0.817|0.183|RT @ericgarland: Trump looks like he swallowed a goldfish and stares at the floor a bit too long.As if maybe a joke has gone too far.
berserk_news||-0.4404|0.182|0.818|0.0|This is what happens when #Donald #Trump attacks a private citizen on Twitter https://t.co/F9CPmeE3Og https://t.co/uiWffpezUb
catlover1943|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
catlover1943|change|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
AberrantEve|TomthunkitsMind|-0.743|0.249|0.671|0.08|RT @TomthunkitsMind: You Can Tell By Trump's Staff Picks That We Are Going To War Within 2 Years. It's A War Cabinet. Get Ready For A Possi
LaEternalSphere|Salon|0.0|0.0|1.0|0.0|RT @Salon: Remember when the anti-globalists were left-wing radicals? https://t.co/eOmlUFsZCb
LaEternalSphere|salon|0.0|0.0|1.0|0.0|RT @Salon: Remember when the anti-globalists were left-wing radicals? https://t.co/eOmlUFsZCb
Truth_of_Truths|realDonaldTrump|0.128|0.108|0.762|0.13|@realDonaldTrump @NBCNightlyNews @CNN there is precisely zero reason to believe anything you say Donald Trump. You'd better resign soon.
SFManeFlame|sarahkendzior|0.0|0.0|1.0|0.0|"RT @sarahkendzior: Two quotes you need to read side by side.1. From Trump 2. From Trump's chief strategist, Steve BannonSpread this wid"
DanielHuculak|SarcasticHoney|0.0|0.0|1.0|0.0|@SarcasticHoney @UniteAlbertans @PC_Alberta and what happened to Mr. Trump in the US he became the president I think
thiswaltz5|quinncy|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
thiswaltz5|palmerreport|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
girishglg|RMConservative|-0.5859|0.178|0.749|0.073|RT @RMConservative: Not all cabinet picks are going 2 b good on every issue. they dont have 2 b. but this one is troubling https://t.co/Rv2
girishglg|t|-0.5859|0.178|0.749|0.073|RT @RMConservative: Not all cabinet picks are going 2 b good on every issue. they dont have 2 b. but this one is troubling https://t.co/Rv2
laysertag|Lrihendry|0.1275|0.113|0.756|0.13|RT @Lrihendry: While shopping 2day I overheard a conv with group saying isn't it great we can say Merry Christmas again &amp; not be afraid! WO
doc_griff_211|comermd|-0.9153|0.444|0.556|0.0|RT @comermd: .@MMFlint plans #DisruptJ20 Trump plans to stop this29 dead &amp; 166 wounded twin bomb attack Istanbul stadium |  https://t.c
doc_griff_211||-0.9153|0.444|0.556|0.0|RT @comermd: .@MMFlint plans #DisruptJ20 Trump plans to stop this29 dead &amp; 166 wounded twin bomb attack Istanbul stadium |  https://t.c
Soitenly125|matthewjdowd|0.4019|0.0|0.886|0.114|"RT @matthewjdowd: Trump calling himself a ""smart person"" reminds me of margaret thatcher: ""if you have to tell people you are a lady, you p"
YellowPup2007|LOLGOP|0.4767|0.0|0.829|0.171|RT @LOLGOP: Ways to get Trump to read intelligence briefs*Centerfolds*Highlights from Hitler speeches*Comment sections*Say they're fro
jlwalker97|VoteHillary2016|0.4019|0.0|0.876|0.124|RT @VoteHillary2016: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.c
jlwalker97||0.4019|0.0|0.876|0.124|RT @VoteHillary2016: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.c
Newyorker2212|ThomJeff7|0.0258|0.09|0.816|0.094|"RT @ThomJeff7: @LionelMedia @YouTube It's over. Bye bye USA. There is no longer objective truth, only spin. Trump (R-Russia) has picked wor"
ValerieEllenLe1|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: GOP Lobbyist requests AG to investigate Trump for political corruption#cnn #msnbc #AMJoy #cnnsotu #thisweek #res
FlyBabyLyn|KeithOlbermann|0.0129|0.08|0.838|0.082|RT @KeithOlbermann: The Russians attacked us to get Trump elected. Here's the evidence @realDonaldTrump is loyal not to us but to them  htt
oufenix|tomtomorrow|-0.7841|0.247|0.703|0.05|RT @tomtomorrow: Thought of what Trump's election means for this country has left me feeling the sort of grief I have felt after death of s
softballscifi|TeaPainUSA|0.5423|0.0|0.769|0.231|"RT @TeaPainUSA: When someone has to tell you they're ""a smart person"", chances are they're not. https://t.co/YPxcAwfAyi"
softballscifi|huffingtonpost|0.5423|0.0|0.769|0.231|"RT @TeaPainUSA: When someone has to tell you they're ""a smart person"", chances are they're not. https://t.co/YPxcAwfAyi"
Jxnewton|kurteichenwald|0.1027|0.133|0.714|0.153|"Oh look, an Australian pol advertising Trump Hotel.No conflicts of interest here. Move on folks.@kurteichenwald https://t.co/zFq3iQOu1C"
Jxnewton|twitter|0.1027|0.133|0.714|0.153|"Oh look, an Australian pol advertising Trump Hotel.No conflicts of interest here. Move on folks.@kurteichenwald https://t.co/zFq3iQOu1C"
richard_lorant|samsteinhp|0.0|0.0|1.0|0.0|"@samsteinhp He knows it. But he also knows that Trump's base will believe it, anyway."
innaroz|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
innaroz|thegatewaypundit|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
_melirubyy_|RUINER|-0.0772|0.075|0.925|0.0|RT @RUINER: When Trump says he's gonna build a wall but you have a trick up your sleeve https://t.co/780ycmYAaJ
_melirubyy_|vine|-0.0772|0.075|0.925|0.0|RT @RUINER: When Trump says he's gonna build a wall but you have a trick up your sleeve https://t.co/780ycmYAaJ
RichardBejah|richardbejah|0.0|0.0|1.0|0.0|#Apple #APPS Apple's Tim Cook among tech executives meeting with Donald Trump on Wedne.. https://t.co/AOvomk74wj https://t.co/ExUpjN6gau
jeffreyrterry|JuddApatow|-0.6486|0.283|0.63|0.087|@JuddApatow This is why Trump won. Most voters can't articulate it but drumbeat of poor policy was hard to miss. https://t.co/Rj54lkYa84
jeffreyrterry|wsj|-0.6486|0.283|0.63|0.087|@JuddApatow This is why Trump won. Most voters can't articulate it but drumbeat of poor policy was hard to miss. https://t.co/Rj54lkYa84
The_Wicker_Man_|InterDD|0.0|0.0|1.0|0.0|@InterDD daqui a pouco ele escreve pro trump querendo dar conselhos de poltica externa pros USA
KauLynn|LadyDoc4Trump|0.0|0.0|1.0|0.0|"RT @LadyDoc4Trump: Our ""president"" says NOTHING, NADA, ZERO about #Christian genocide by his Muslim brothers.#Trump speaks #Truth on it."
NicolasRobidoux|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
anesam98|NicholsUprising|-0.296|0.115|0.885|0.0|RT @NicholsUprising: And it was a union leader from Indiana who dared to say the emperor has no clothes...https://t.co/Lx3wWj4rCc
anesam98|thenation|-0.296|0.115|0.885|0.0|RT @NicholsUprising: And it was a union leader from Indiana who dared to say the emperor has no clothes...https://t.co/Lx3wWj4rCc
slidewinding|JYSexton|0.5106|0.0|0.883|0.117|RT @JYSexton: It's not even a mystery how Trump was able to finally break the tether of trust between his voters and the media. It was beyo
MikeMongo|andyoutis|0.0|0.0|1.0|0.0|"RT @andyoutis: If you have 7 min, this thread on what led to the election of Trump, Russia's likely strategy, and where we go from here is"
Kenshiro73|JSavoly|-0.0258|0.114|0.778|0.108|RT @JSavoly: Top Republicans Just Demanded An Investigation Into Russia's Pro-Trump Interference #StollenElection #ComradeTrump  https://t.
Kenshiro73||-0.0258|0.114|0.778|0.108|RT @JSavoly: Top Republicans Just Demanded An Investigation Into Russia's Pro-Trump Interference #StollenElection #ComradeTrump  https://t.
tyme11|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
tyme11||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
crichlow|liamstack|0.0772|0.105|0.739|0.156|RT @liamstack: Now that Twitter has cracked down on the pro-Trump bots the top replies to @realDonaldTrump are mostly comedians mocking him
dremtee|toralvaria|0.7003|0.0|0.721|0.279|"RT @toralvaria: Trump is changing and writing new rules, declines receiving daily intelligence briefings. Interesting actually.  https://t."
dremtee||0.7003|0.0|0.721|0.279|"RT @toralvaria: Trump is changing and writing new rules, declines receiving daily intelligence briefings. Interesting actually.  https://t."
k_r_eckert|chavezglen1755|0.2103|0.0|0.831|0.169|RT @chavezglen1755: WHY VLADIMIR PUTINS RUSSIA IS BACKING DONALD TRUMPhttps://t.co/FkSdXjOmCg
Tamaraciocci|melreynoldsU|-0.5423|0.143|0.857|0.0|"RT @melreynoldsU: Rubio, McCain and Graham are not up for reelection, they literally could destroy Donald Trump's time in the White House a"
cthulhucloaca|cushbomb|-0.5267|0.159|0.841|0.0|@cushbomb we need a conspiracy theory saying the FSB controls Trump because Melania was a matahari who turned him into a Krok-head
Monte_Alto|realDonaldTrump|-0.4404|0.225|0.775|0.0|#Trump's Dirty money: @realDonaldTrump and the Kazakh connection https://t.co/BQ4NRpeGlv via @FT
Monte_Alto|ft|-0.4404|0.225|0.775|0.0|#Trump's Dirty money: @realDonaldTrump and the Kazakh connection https://t.co/BQ4NRpeGlv via @FT
LegendaryClan__|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
boy45691713|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
boys59483916|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
NOMADD11|NOMADD11|0.0|0.0|1.0|0.0|@NOMADD11 @maddow @NYTupelo7 @morgfair @samsteinhp @BBCWorld @Elise_Jordan @cristina5411 @SHAQ @chrislhayes: TRUMP SECRET PLANS 4 AMERICANS!
mtighe15|ezlusztig|-0.6249|0.17|0.83|0.0|"RT @ezlusztig: Purely on the basis of information publicly available - just the tip of an iceberg, presumably - Obama could devastate Trump"
rachel1970|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
V_of_Europe|thegatewaypundit|-0.0772|0.279|0.508|0.213|Trump: Democrats Just Suffered One of Greatest Defeats in History of Politics  https://t.co/L255CE0Kjp
Burger_Buzz|Cernovich|0.128|0.0|0.842|0.158|"@Cernovich Trump is a Russian agent. Tread carefully, Trump Traitors."
cjedwards65|kurteichenwald|-0.128|0.181|0.7|0.119|RT @kurteichenwald: The intel briefings include critical information designed to keep our troops safe. It changes every day. Trump ignores
ahernandez85a|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
ahernandez85a|thegatewaypundit|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
MESoundX4|AnaRent|0.0|0.0|1.0|0.0|RT @AnaRent: Hay esperanza! @washingtonpost revela que la #CIA encontr que #Rusia intervino en las Elecciones de #EU para favorecer a Don
EnriqueM77|TheMarkRomano|0.2263|0.087|0.786|0.127|"RT @TheMarkRomano: NBC news still pushing the ""Trump supporters are Klan members and White supremacists"" propaganda.NBC, you guys are dis"
IsaLeeWolf|riotwomennn|0.5622|0.0|0.846|0.154|"RT @riotwomennn: Retweet &amp; post on your social media.  This is EASY.  Takes 5 minutes.  Go to https://t.co/DoLmGiiYVf  Fill this out, hit s"
IsaLeeWolf|asktheelectors|0.5622|0.0|0.846|0.154|"RT @riotwomennn: Retweet &amp; post on your social media.  This is EASY.  Takes 5 minutes.  Go to https://t.co/DoLmGiiYVf  Fill this out, hit s"
DtRh321|textifyer59|0.0|0.0|1.0|0.0|"@textifyer59 @LouiseMensch ""secret"" trump server? otherwise known as server."
GregPoliteia|RoseAnnDeMoro|0.2023|0.0|0.899|0.101|"RT @RoseAnnDeMoro: For someone who wants to #draintheswamp, Trump keeps reaching into Goldman Sachs for appointments: https://t.co/UQwySYRC"
GregPoliteia|t|0.2023|0.0|0.899|0.101|"RT @RoseAnnDeMoro: For someone who wants to #draintheswamp, Trump keeps reaching into Goldman Sachs for appointments: https://t.co/UQwySYRC"
JacobDanielsOR|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
LaVerneWright13|Worldofcraze|0.3818|0.0|0.885|0.115|RT @Worldofcraze: Trump locking every job in the government to ensure full control to achieve all his goals unchallenged and unpunished.T
TimothyKopp2|JrcheneyJohn|0.0|0.0|1.0|0.0|RT @JrcheneyJohn: The #FakeNews Media has been Neutered by Trump and they have become Irrelevant #TrumpEffect  https://t.co/8ArN8MrraK
TimothyKopp2|twitter|0.0|0.0|1.0|0.0|RT @JrcheneyJohn: The #FakeNews Media has been Neutered by Trump and they have become Irrelevant #TrumpEffect  https://t.co/8ArN8MrraK
Piter432YT|TygodnikLisicki|0.0|0.0|1.0|0.0|RT @TygodnikLisicki: TYLKO W DO RZECZY Matthew Tyrmand rozmawia z Donald J. Trump o Polsce: Bardzo przychylnie wypowiada si o... https
iu70us|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
iu70us|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
MonicaFitz1|BelkissObadia|-0.4588|0.125|0.875|0.0|RT @BelkissObadia: #TRUMPLEAKS Donald Trump will be the reason our country is going to get attacked because of his narcissistic madman beha
HonkyTonkNights|breitbart|0.7579|0.0|0.629|0.371|Conway: Conclusion Russia Was Acting to Help Trump Win Election Are 'Ridiculous' https://t.co/5D0oemzu2I
vtti|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
vtti|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
luishlear|jimpavia|0.0|0.0|1.0|0.0|"RT @jimpavia: Trump says Wall Street Journal doesn't ""understand business"" https://t.co/Au9HPkKf5D"
luishlear|cnbc|0.0|0.0|1.0|0.0|"RT @jimpavia: Trump says Wall Street Journal doesn't ""understand business"" https://t.co/Au9HPkKf5D"
paintbygretzky|StacyLeMelle|0.0|0.0|1.0|0.0|RT @StacyLeMelle: THIS IS WHAT I'M TALKING ABOUT! @VanJones68 Bravo!! @TheChrisSuprun #hamiltonelectors #ElectoralCollege https://t.co/Wh
paintbygretzky|t|0.0|0.0|1.0|0.0|RT @StacyLeMelle: THIS IS WHAT I'M TALKING ABOUT! @VanJones68 Bravo!! @TheChrisSuprun #hamiltonelectors #ElectoralCollege https://t.co/Wh
Frannn_____|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
rafacapozzi|labanda|-0.4184|0.148|0.852|0.0|Yo no se que es peor que ganar trump o que @labanda fuera un desastre como esta!! ASCOOOOO
KayHillYes|HamiltonElector|-0.296|0.099|0.901|0.0|RT @HamiltonElector: We've crossed the threshold. There is no going back. Trump must never become POTUS. RT to let #hamiltonelectors know y
cosmokramerss|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
catheri81371820|Trollin_Trump|-0.6705|0.251|0.643|0.106|"@Trollin_Trump The worst thing you can do to a narcissist is make fun of them .They hate it ,it fracture there ego.Keep it coming."
ErrantStrategry|jayrosen_nyu|-0.2144|0.074|0.926|0.0|"RT @jayrosen_nyu: 19/ The problem is not at the level ""how to cover Trump,"" but how to recover conditions in which anything journalists do"
MargoErickson9|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Sam777rt|DanScavino|0.5106|0.163|0.555|0.282|"RT @DanScavino: ""NO DREAM is too big, NO CHALLENGE is too great. Nothing we want for our future is BEYOND OUR REACH."" Donald J. Trump, Pre"
DRocks777|SarahLerner|0.0|0.0|1.0|0.0|"RT @SarahLerner: So to recap, Russia intervened in our election to achieve a specific outcome: Elect Donald Trump. How are people not more"
DonnieBolena|foxnews|-0.1511|0.104|0.825|0.071|The media exaggerates everything they say!GOP senators challenge Trump on secretary of state prospect's Russia ties. https://t.co/nsjldSkQYi
SmokinSam420|TrumpNewMedia|-0.6833|0.236|0.764|0.0|RT @TrumpNewMedia: 3 #Traitors @SenJohnMcCain @LindsayGrahamSC @marcorubio WARS cost #America $6 Trillion dollars! #Reuters #GOP #Trump #MA
ArtsLetter|thedailybeast|-0.7096|0.396|0.604|0.0|RT @thedailybeast: Carl Bernstein: Trump's lies worse than Nixon's:  https://t.co/wBaRkFjidX https://t.co/8lgakwPLpe
ArtsLetter|thedailybeast|-0.7096|0.396|0.604|0.0|RT @thedailybeast: Carl Bernstein: Trump's lies worse than Nixon's:  https://t.co/wBaRkFjidX https://t.co/8lgakwPLpe
mzzcocoa|netw3rk|-0.4215|0.304|0.543|0.152|RT @netw3rk: 2016Media: white supremacists dress nice nowTeen Vogue: Trump is destroying democracy
millerjr99|nbcnews|-0.8237|0.353|0.647|0.0|You can't make this shit up!!! #trumpgretsTrump (Wrongly) Criticized Obama for Not Attending Intel Briefings - https://t.co/4f3fRXeaNm
EchoPapaDelta|DRUDGE_REPORT|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: SPY GAMES https://t.co/Hjpfjm4G5M
EchoPapaDelta|cnn|0.0|0.0|1.0|0.0|RT @DRUDGE_REPORT: SPY GAMES https://t.co/Hjpfjm4G5M
Teeda100|tonyschwartz|-0.296|0.091|0.909|0.0|RT @tonyschwartz: I don't believe anything Donald Trump says. Not one word. It is all manipulation and mind games all the time. (Same for K
nmclaughlin04|phillydotcom|0.0|0.0|1.0|0.0|"Trump, Putin, McConnell and the plot against America https://t.co/pOTt9Nhrcy via @phillydotcom"
nmclaughlin04|philly|0.0|0.0|1.0|0.0|"Trump, Putin, McConnell and the plot against America https://t.co/pOTt9Nhrcy via @phillydotcom"
SummerCampus_|bloomberg|-0.34|0.179|0.821|0.0|business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/WQtS9dzzvk https://t.co/Atwcgt1muR
Cobra1A|mormorlady|-0.6542|0.235|0.687|0.078|@mormorlady @MikeCarlton01 He is now in heaven since  Trump  became President   ..the man is brain dead but Turnbull  is scared of him
SlyDurin|kurteichenwald|0.126|0.146|0.687|0.167|"RT @kurteichenwald: Putin staff consultant re: Trump choices: ""This is a fantastic team!""Remember when Romney said Russia biggest threat?"
katherinejnowak|teeg_dougland|-0.8126|0.381|0.619|0.0|"@teeg_dougland @neeratanden 45. highlighting trump's strengthsunpredictable, bad boy, etcas any kind of character assassination"
WendyBrandes|summerbrennan|-0.5277|0.206|0.726|0.069|RT @summerbrennan: This isn't good. Not at all: Russia tests new underwater nuclear drone amid growing tensions with the West https://t.co/
WendyBrandes|t|-0.5277|0.206|0.726|0.069|RT @summerbrennan: This isn't good. Not at all: Russia tests new underwater nuclear drone amid growing tensions with the West https://t.co/
WendyBrandes|JRubinBlogger|-0.0516|0.216|0.632|0.153|RT @JRubinBlogger: Trump's Disregard of Intel Findings is 'Extraordinarily Beneficial to Russian Propaganda' https://t.co/vh8V5xWdH1 Schiff
WendyBrandes|mediaite|-0.0516|0.216|0.632|0.153|RT @JRubinBlogger: Trump's Disregard of Intel Findings is 'Extraordinarily Beneficial to Russian Propaganda' https://t.co/vh8V5xWdH1 Schiff
SarahGBloom|SalAntoni0|-0.0572|0.08|0.92|0.0|RT @SalAntoni0: The side of Donald Trump the media doesn't want you to see  https://t.co/Yvd3EhetEF
SarahGBloom|twitter|-0.0572|0.08|0.92|0.0|RT @SalAntoni0: The side of Donald Trump the media doesn't want you to see  https://t.co/Yvd3EhetEF
RealKin88|haydenblack|0.7184|0.0|0.731|0.269|"RT @haydenblack: #Trump now tweeting that the CIA is ""highly overrated"" and should apologize to Russia which should be a ""safe and special"
NicholasMe|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
HGTomato|liamstack|0.0772|0.105|0.739|0.156|RT @liamstack: Now that Twitter has cracked down on the pro-Trump bots the top replies to @realDonaldTrump are mostly comedians mocking him
rhetoricAli|MichaelSkolnik|-0.4588|0.125|0.875|0.0|RT @MichaelSkolnik: Many Republicans are going to have a rude awakening when they finally realize what we all have known. Trump is putting
NastyBoof1970|GovHowardDean|0.0|0.0|1.0|0.0|RT @GovHowardDean: Why Putin Prefers Trump https://t.co/U2B9kZg38D
NastyBoof1970|politico|0.0|0.0|1.0|0.0|RT @GovHowardDean: Why Putin Prefers Trump https://t.co/U2B9kZg38D
mishayah|Lagartija_Nix|-0.4767|0.181|0.819|0.0|RT @Lagartija_Nix: Trump Blasts CNN for Fake News Report on The Apprentice https://t.co/OZtYVtbXvn via @LifeZette
mishayah|lifezette|-0.4767|0.181|0.819|0.0|RT @Lagartija_Nix: Trump Blasts CNN for Fake News Report on The Apprentice https://t.co/OZtYVtbXvn via @LifeZette
Dhriyamana|mitchellvii|-0.7351|0.22|0.78|0.0|RT @mitchellvii: I don't get it.  The Media is using the same attacks against Trump that failed during the election.  They need to hire bet
jackhenrynola|quinncy|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
jackhenrynola|palmerreport|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
bhavesh1968p|ckmarie|0.6892|0.0|0.562|0.438|@ckmarie @JoyAnnReid that trump is awesome !!
binamutha|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
S29Allen|rudepundit|-0.765|0.248|0.752|0.0|"RT @rudepundit: Maybe Trump is too dumb to understand that the word ""intelligence"" isn't meant as an insult to those being briefed."
LatorreNina|NathanZed|0.0|0.0|1.0|0.0|RT @NathanZed: Trump really out here having meetings with four Lex Luthor's https://t.co/7vbYrU6eSB
LatorreNina|twitter|0.0|0.0|1.0|0.0|RT @NathanZed: Trump really out here having meetings with four Lex Luthor's https://t.co/7vbYrU6eSB
cagneylou|alternet|-0.4215|0.149|0.851|0.0|5 Ways Hillary Clinton Can Mock Thin-Skinned Trump to Make Him Go Bonkers at Tonight's Debate @alternet https://t.co/PueNYJEYij
cagneylou|alternet|-0.4215|0.149|0.851|0.0|5 Ways Hillary Clinton Can Mock Thin-Skinned Trump to Make Him Go Bonkers at Tonight's Debate @alternet https://t.co/PueNYJEYij
FosterF31757930|LouDobbs|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
FosterF31757930|theconservativetreehouse|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
trishmaximum|Reuters|0.2023|0.0|0.878|0.122|RT @Reuters: Top tech executives to attend Trump summit on Wednesday: Recode https://t.co/nhMs2ST41h https://t.co/pEFtYNUBVL
trishmaximum|reuters|0.2023|0.0|0.878|0.122|RT @Reuters: Top tech executives to attend Trump summit on Wednesday: Recode https://t.co/nhMs2ST41h https://t.co/pEFtYNUBVL
SusanCarver19|Amplitude350Lee|-0.4767|0.129|0.871|0.0|RT @Amplitude350Lee: @AirborneChick @bsbafflesbrains  How anyone could watch what Trump has done and still say HRC is worse is beyond my co
noisyparker|chrisantenucci|0.2023|0.0|0.909|0.091|RT @chrisantenucci: https://t.co/TnJqh2ZavIThis is an important article for anyone who wants to understand why our intel agencies have be
noisyparker|t|0.2023|0.0|0.909|0.091|RT @chrisantenucci: https://t.co/TnJqh2ZavIThis is an important article for anyone who wants to understand why our intel agencies have be
mtada71|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
MrCoolcasi|factcheckdotorg|-0.5859|0.194|0.806|0.0|RT @factcheckdotorg: Trump again doubted that Russia was behind the hacked emails during the election. Here's the evidence that it was: htt
outerspacemanII|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
RWonder777|fxn.ws|-0.5267|0.173|0.827|0.0|Trump filling his Cabinet with ObamaCare foes @fxn.ws - Obamacare needs to be changed. Cost too steep for middle class &amp; taxpayers to pay.
betsyanne|latimes|0.0|0.0|1.0|0.0|"'A dog and pony show,' lawyer in class-action suit says, recalling Trump University seminar https://t.co/sV1GABzqsl"
EmmeWinch|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
EmmeWinch||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
Daniel7964|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
Sp3ck_Sec|t|0.0|0.0|1.0|0.0|"CIA report: Russia helped Trump in Presidential election: https://t.co/HXpQhQW04JA month later result of US Presidential election, Ameri"
manish_vij|HeerJeet|0.7003|0.0|0.707|0.293|"RT @HeerJeet: Well, at least the Russians are happy with Tillerson's (possible) appointment    : Trump continues to a"
Bellalindafox|dolceamori|-0.6597|0.265|0.735|0.0|RT @dolceamori: Troubling op-ed in Trump in-laws newspaper calls for FBI crackdown on anti-Trump protests https://t.co/n7Ny9b0ci5 #Resist
Bellalindafox|rawstory|-0.6597|0.265|0.735|0.0|RT @dolceamori: Troubling op-ed in Trump in-laws newspaper calls for FBI crackdown on anti-Trump protests https://t.co/n7Ny9b0ci5 #Resist
raemadema|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
readbetsyread|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
swissifg|marketwatch|-0.0258|0.14|0.725|0.135|Trump is inspiring investors to abandon the post-financial-crisis search for yield and cycling into big bets: https://t.co/dmcUEQ7k8I
LyraSona|asamjulian|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
LyraSona|twitter|0.1779|0.098|0.765|0.137|"RT @asamjulian: Russophobia is actually a form of xenophobia, something liberals like to accuse Trump of. https://t.co/RWFlg7Lx97"
bibi4Trump|insider|0.0|0.0|1.0|0.0|https://t.co/AiKIM4w25x
LisaMoraitis1|HamiltonElector|0.2298|0.123|0.757|0.12|"RT @HamiltonElector: Mr. Trump you are hardly a genius, no matter what Comrade Putin says.  We are smarter than you. We are #hamiltonelecto"
mimizelman|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
MichaelBarlow42|nytimesbusiness|0.4019|0.0|0.886|0.114|"RT @nytimesbusiness: CEOs see a Field of Dreams economy under Trump. If you are a Republican, this is the beginning of a golden age. http"
andykhouri|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
andykhouri||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
elysium55|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
LauraDuet1|KaraCalavera|0.3182|0.0|0.887|0.113|"RT @KaraCalavera: I'm sure they also called for an investigation into Trump's business dealings. Oh, they didn't? Hmm... https://t.co/W3q"
LauraDuet1|t|0.3182|0.0|0.887|0.113|"RT @KaraCalavera: I'm sure they also called for an investigation into Trump's business dealings. Oh, they didn't? Hmm... https://t.co/W3q"
AndreaDBergman|kurteichenwald|0.4215|0.0|0.877|0.123|RT @kurteichenwald: .@SenJohnMcCain - briefed on intel - say on air that he knows evidence of Russian interference and its true. Trump team
Lisa_Iannucci|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
ggprez|TayTay78730804|0.4084|0.104|0.702|0.195|RT @TayTay78730804: #SundayMorning I find it funny how liberals cry about trump wanting to build a wall. It's OK for them to put one up tho
eprophotog|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: US Senators letter to Senate leaders-investigate Trump for Russian espionage#cnn #msnbc #AMJoy #cnnsotu #thiswee
Inked1BNA|hollyoptix|-0.4404|0.255|0.607|0.138|RT @hollyoptix: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/4J4gQ
Inked1BNA|t|-0.4404|0.255|0.607|0.138|RT @hollyoptix: US Justice Department: Prosecute Trump for illegal activities before the Dec. 19 Electoral College Vo... https://t.co/4J4gQ
ArgentinaPatito|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
CIMAGES|AP|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
CIMAGES|t|-0.4939|0.151|0.849|0.0|"RT @AP: #AP10Things: Trump rejects intel, lawmakers vow probe of Russia hacking; IS militants retake ancient Syrian city. https://t.co/3NQ7"
AJ_Rutten|ErinSchrode|0.4342|0.154|0.557|0.289|"RT @ErinSchrode: THIS. IS. TERRIFYING. Trump will NOT receive daily intelligence briefings bc You know, Im, like, a smart person."" https"
Royce_Yoho|kurteichenwald|-0.5423|0.176|0.824|0.0|"RT @kurteichenwald: Fox/Cheney went nuts when found out Obama got intel briefings in writing, rather than read to him. But Trump no briefin"
orlandolatino|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Anyone else unnerved by all the tech CEOs making the pilgrimage to Trump Tower?
ggbootsrock|LouDobbs|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
ggbootsrock|theconservativetreehouse|0.3612|0.0|0.872|0.128|RT @LouDobbs: The Natural - President Donald Trump TV Appearance at Army -vs- Navy Game https://t.co/sSg1mCoWfb via @thelastrefuge2 #MAGA @
bdanaher17|reuters|0.2732|0.0|0.811|0.189|Rick Perry a leading candidate for U.S. energy post: source https://t.co/12cgLGV6Ft
MrJamesJoint|nbcsnl|0.4588|0.0|0.769|0.231|"RT @nbcsnl: Welcome to the Trump administration, Walter White. #CenaOnSNL https://t.co/aPaceUQcO0"
MrJamesJoint|twitter|0.4588|0.0|0.769|0.231|"RT @nbcsnl: Welcome to the Trump administration, Walter White. #CenaOnSNL https://t.co/aPaceUQcO0"
RightSideFTW|JayJ2Great|0.7452|0.0|0.784|0.216|@JayJ2Great @CP24 Trump loves Canada and isnt to be feared - took old C PM's to get that sorted.  Now we need a PM to work with him
layna_bayna|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
layna_bayna||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
alecrider|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
alecrider||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
MRICTPET|AAPsyc|0.8374|0.114|0.504|0.381|@AAPsyc don't you understand? Your degree of unhappiness is proportional to my degree of happiness LOL love my trump...
PSemec|ScottCPhilips|0.0|0.0|1.0|0.0|"@ScottCPhilips @AlecMacGillis The media gave Trump SO MUCH coverage of each of his ""missteps"", ppl were desensitized: he wrote off almost"
cclement873|vivelafra|-0.6486|0.194|0.806|0.0|"RT @vivelafra: BIG 6: After criminally colluding with his opponent for 18 months, MSM is now trying to suggest #Trump had an unfair advanta"
JimJinksCT|twitter|-0.6249|0.316|0.563|0.122|Good headline but undersells the misery embodied by Trump. #Trumpocalyp https://t.co/IGWHt2VD5l
FOX61News|fox61|0.0|0.0|1.0|0.0|Trump: 'Nobody really knows' if climate change is real https://t.co/Kjt8Lpyxw5 https://t.co/SW18wXQGq6
dbart59|_Makada_|-0.296|0.115|0.826|0.06|"RT @_Makada_: President-Elect Trump: It's ridiculous to say Russia intervened in the election, I think it's just another excuse. We had a m"
pisannd5|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
beemerjean|whattrumpdid|0.0772|0.137|0.711|0.152|RT @whattrumpdid: Our #delusionistinchief has a bit of an ego problem https://t.co/Ol3jKVnXCm welcome to #TrumpNation #thenewswamp #theresi
beemerjean|huffingtonpost|0.0772|0.137|0.711|0.152|RT @whattrumpdid: Our #delusionistinchief has a bit of an ego problem https://t.co/Ol3jKVnXCm welcome to #TrumpNation #thenewswamp #theresi
thinkerdamous|cnn|-0.5356|0.219|0.687|0.094|What would a real leader do? Not Trump https://t.co/VyMFn0d7H1 Trump is an incredibly stupid &amp; naive person. Leaders 1st job is to protect.
MLorance|kurteichenwald|0.5574|0.0|0.847|0.153|"RT @kurteichenwald: If Trump started getting praise 4  appointments from ISIS, do you think Fox News would start running stories about how"
katriord|ericgarland|-0.2052|0.114|0.805|0.08|"RT @ericgarland: And now, it's December 11th. Trump says he don't need no stinkin' intel agencies. Russia (BWA HAHAHAHAAAA) blames Ukrain"
Patar4950|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
supercub666|johncheese|-0.8625|0.336|0.664|0.0|"RT @johncheese: If Stephen Hawking told Trump he's wrong about black holes, Trump would call him an idiot. ""He's anti-science. A moron. Big"
JbthomJohn|demandprogress|-0.3595|0.142|0.858|0.0|Sign now: Tell tech companies to refuse to build Trump's Muslim registry! https://t.co/2n3CfYr00A via @demandprogress #NoMuslimRegistry
JbthomJohn|act|-0.3595|0.142|0.858|0.0|Sign now: Tell tech companies to refuse to build Trump's Muslim registry! https://t.co/2n3CfYr00A via @demandprogress #NoMuslimRegistry
lauraannmariee|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
Phillipdrphl|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
ColBannister|realJeffreyLord|-0.0387|0.183|0.678|0.139|@realJeffreyLord @Mediaite but you are the one thing I miss on @cnn Jeff- you are a true professional &amp; fought for President-Elect Trump
Sbecher|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
TrdngDrivatives|EnviroNews|0.4215|0.098|0.684|0.218|RT @EnviroNews: #Trump Portfolio Riddled w/ Oil Stocks - Conflict of Interest for Him to Sign Energy Bills? https://t.co/jKKyuJOZaT https:/
TrdngDrivatives|environews|0.4215|0.098|0.684|0.218|RT @EnviroNews: #Trump Portfolio Riddled w/ Oil Stocks - Conflict of Interest for Him to Sign Energy Bills? https://t.co/jKKyuJOZaT https:/
bradpotterbaum|reddit|0.296|0.0|0.845|0.155|Elon Musk To Join Trumps Tech-Industry Summit In New York This Week https://t.co/rdZ75dO3mU
nakedlaughing|laurine3215|-0.7213|0.267|0.668|0.065|"RT @laurine3215: Sad that even Trump supporters REALLY don't believe him, but don't want to look stupid for voting for him.That is why they"
slowbuck|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
michaelob123|pixelatedboat|-0.4585|0.167|0.833|0.0|RT @pixelatedboat: I read the 12th Amendment and technically neither Clinton nor Trump won the election: https://t.co/fKieKK3fEH
michaelob123|twitter|-0.4585|0.167|0.833|0.0|RT @pixelatedboat: I read the 12th Amendment and technically neither Clinton nor Trump won the election: https://t.co/fKieKK3fEH
JudyHistorian|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
JudyHistorian|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
srekita7|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
KathyLittle18|WG_Burton|0.1531|0.0|0.833|0.167|RT @WG_Burton: A Carefully Planned Operation to Prevent President-elect Donald Trumps Accession to the White House?https://t.co/HQHpFUBoH
KathyLittle18|t|0.1531|0.0|0.833|0.167|RT @WG_Burton: A Carefully Planned Operation to Prevent President-elect Donald Trumps Accession to the White House?https://t.co/HQHpFUBoH
vasiliy_b|Bernies4_Trump|0.0|0.0|1.0|0.0|@Bernies4_Trump @EcuadorDeb @MissLizzyNJ the crucial point -- it were Russian servicemen.
Aroberts521|washingtonpost|0.8481|0.0|0.62|0.38|If only modern politician had the courage to avail themselves the system our founding fathers brilliantly created. https://t.co/CRoRX2J984
Patkrick|Salon|0.0|0.0|1.0|0.0|@Salon Trump President Nahhhhh!!!!
OrmondDerrick|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
LIVEdude|yahoo|0.4019|0.0|0.87|0.13|Stay sharp out there. The #FED may pop some balloons on their way through the party. #InterestHike #PartyIsOverParty https://t.co/SPKL5uSwMR
Shelleypg19|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Shelleypg19||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
jknizer|lbo-news|0.0|0.0|1.0|0.0|https://t.co/AVuEHvu6kA
dolceamori|occupydemocrats|0.25|0.079|0.787|0.135|FOX Just Called Out Trump For His Pay For Play Hypocrisy To His Face - https://t.co/MxKWQpMQrO  #Resist
DAILYBLUEblog|RalfThePowerful|-0.2023|0.083|0.917|0.0|"RT @RalfThePowerful: When confronted with evidence that Russia worked to elect him, rather than ""I can't be bought,"" Trump's statement was"
AlwaystrumpOrg|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
longshipdriver|Jodzio|-0.8625|0.346|0.654|0.0|"RT @Jodzio: Putin must have 'smoking gun"" that can ruin Trump. Probably sex related. But worse than anything that has been exposed so far."
pufftrishy|aravosis|0.4767|0.0|0.846|0.154|RT @aravosis: Kellyanne Conway says Trump is going to put his own people in the intelligence community https://t.co/3wew3gUmr7
pufftrishy|shareblue|0.4767|0.0|0.846|0.154|RT @aravosis: Kellyanne Conway says Trump is going to put his own people in the intelligence community https://t.co/3wew3gUmr7
LozierJeannine|AriMelber|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
LozierJeannine|t|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
sherrilee7|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
BSAFunds|marketwatch|-0.0258|0.14|0.725|0.135|Trump is inspiring investors to abandon the post-financial-crisis search for yield and cycling into big bets: https://t.co/Pghv5mpIHD M
CJThompson87|marklevinshow|-0.6369|0.276|0.724|0.0|RT @marklevinshow: More Goldman Sachs appointments; I thought Trump hated Goldman Sachs https://t.co/d93fhyI6cG
CJThompson87|conservativereview|-0.6369|0.276|0.724|0.0|RT @marklevinshow: More Goldman Sachs appointments; I thought Trump hated Goldman Sachs https://t.co/d93fhyI6cG
carolina_brenna|CDoranHarader|-0.946|0.571|0.429|0.0|RT @CDoranHarader: Muslim extremist who lied about hate crime goes into hiding to avoid being arrested for hoax... https://t.co/dH4eItOt4B
carolina_brenna|linkis|-0.946|0.571|0.429|0.0|RT @CDoranHarader: Muslim extremist who lied about hate crime goes into hiding to avoid being arrested for hoax... https://t.co/dH4eItOt4B
incrementable|markmobility|0.3818|0.0|0.874|0.126|"RT @markmobility: While Trump promises to bring jobs home, he quietly hires 64 foreign workers at Mar-a-Lago https://t.co/2IpSahqgBW https:"
incrementable|mypalmbeachpost|0.3818|0.0|0.874|0.126|"RT @markmobility: While Trump promises to bring jobs home, he quietly hires 64 foreign workers at Mar-a-Lago https://t.co/2IpSahqgBW https:"
macmcd|DailyNewsBin|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
macmcd|palmerreport|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
charmingred|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
YvetteKopp|moderatemama|0.5719|0.0|0.748|0.252|@moderatemama have you watched this video from Russia after Trump won? https://t.co/tdxv2h3NNk
YvetteKopp|youtube|0.5719|0.0|0.748|0.252|@moderatemama have you watched this video from Russia after Trump won? https://t.co/tdxv2h3NNk
ANUR01|huffingtonpost|0.0|0.0|1.0|0.0|https://t.co/dfqiISXKdO
RobertA87413263|realjunsonchan|-0.4215|0.272|0.545|0.183|RT @realjunsonchan: Brave man Joe Scarborough risks his own life to tell truth against feral idiot fake news media. #Trump #maga #underdoge
CR710349|France4Hillary|0.4753|0.0|0.86|0.14|RT @France4Hillary: BREAKING: #Hillary's popular vote lead over Trump is now close to 3 million votes! #HillaryWon - SHE'S THE PEOPLE'S CHO
totoqro|actualidad|0.0|0.0|1.0|0.0|https://t.co/CFnUzHd18M
Girl__III|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Girl__III||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
ribcagestyles|glennspizza|-0.1027|0.167|0.833|0.0|"RT @glennspizza: ""maggie for president"" trump is shook"
DinaJon60818043|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
DinaJon60818043|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
RyanResign|TrumpNewMedia|-0.6833|0.236|0.764|0.0|RT @TrumpNewMedia: 3 #Traitors @SenJohnMcCain @LindsayGrahamSC @marcorubio WARS cost #America $6 Trillion dollars! #Reuters #GOP #Trump #MA
Tuna_Ghost|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Alehandro9390|Magiq1|-0.296|0.206|0.688|0.106|"RT @Magiq1: What time is it. @Magiq1 Abortion Foes, Emboldened by Trump, Promise Onslaught of Tough Restrictions https://t.co/JtORjbW2Ap"
Alehandro9390|nytimes|-0.296|0.206|0.688|0.106|"RT @Magiq1: What time is it. @Magiq1 Abortion Foes, Emboldened by Trump, Promise Onslaught of Tough Restrictions https://t.co/JtORjbW2Ap"
JPegios|LDrogen|0.7096|0.0|0.731|0.269|RT @LDrogen: Good luck to the coal miners who got conned by Trump Fully autonomous coal mine https://t.co/g7QXQH3jY5
JPegios|twitter|0.7096|0.0|0.731|0.269|RT @LDrogen: Good luck to the coal miners who got conned by Trump Fully autonomous coal mine https://t.co/g7QXQH3jY5
PattiPropst|lifezette|0.0|0.0|1.0|0.0|https://t.co/2QEOgmKmGn
ekingc|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
ekingc|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
MiaShaw|oliverdarcy|0.0|0.0|1.0|0.0|RT @oliverdarcy: Rubio chides Trump for boasting about likely sec of state pick's relationship with Putin https://t.co/XkPiqeBDro
MiaShaw|businessinsider|0.0|0.0|1.0|0.0|RT @oliverdarcy: Rubio chides Trump for boasting about likely sec of state pick's relationship with Putin https://t.co/XkPiqeBDro
FrancesRauer|HamiltonElector|-0.4401|0.115|0.843|0.042|RT @HamiltonElector: RT The only thing that matters now is educating EVERYONE that Donald Trump is not President yet. He has not won. #Dec1
SandraW11075083|funder|-0.3237|0.109|0.891|0.0|RT @funder: #TRUMPLEAKS EXPOSED THIS! Carrier Got Taxpayer Handout Because Trump Owns Stock In Their Parent Company #cnn #msnbc https://t.c
SandraW11075083||-0.3237|0.109|0.891|0.0|RT @funder: #TRUMPLEAKS EXPOSED THIS! Carrier Got Taxpayer Handout Because Trump Owns Stock In Their Parent Company #cnn #msnbc https://t.c
DivaDollar|HuffPostPol|0.0|0.0|1.0|0.0|"RT @HuffPostPol: Trump says ""nobody really knows"" if climate change is real (It is.) https://t.co/zstqb4f01i https://t.co/nQg5iMdLXx"
DivaDollar|m|0.0|0.0|1.0|0.0|"RT @HuffPostPol: Trump says ""nobody really knows"" if climate change is real (It is.) https://t.co/zstqb4f01i https://t.co/nQg5iMdLXx"
svenosaurus|twitter|0.8814|0.0|0.624|0.376|"Emcee Trump: Audience thinks T Rex is too close to my friend Putin? OK, then the winner is John Bedlam! https://t.co/Dk0FosUPMY"
kals55|NPR|-0.1779|0.124|0.876|0.0|"RT @NPR: As Trump Dismisses CIA, Congress Looks To Confront Russian Cyberattacks https://t.co/CLExlZVvHT"
kals55|npr|-0.1779|0.124|0.876|0.0|"RT @NPR: As Trump Dismisses CIA, Congress Looks To Confront Russian Cyberattacks https://t.co/CLExlZVvHT"
ElisaPerezG1|PressTV|0.4939|0.0|0.775|0.225|@PressTV Trump can be 'its only one friend' or 'its imaginary friend'.
facklernyt|ftasia|0.34|0.0|0.882|0.118|"RT @ftasia: Trump puts four-decade old ""One China"" policy in play: Trumps position is you can trade anything  https://t.co/5LQEN0Pjmy"
facklernyt|ft|0.34|0.0|0.882|0.118|"RT @ftasia: Trump puts four-decade old ""One China"" policy in play: Trumps position is you can trade anything  https://t.co/5LQEN0Pjmy"
jhrusher|Politics_PR|0.0|0.0|1.0|0.0|@Politics_PR recounts really? at who's request are the counts being done? steins or clinton? and trump isn't afraid of them so answer
Pink22Karen|rdlaing|-0.8271|0.34|0.584|0.076|"RT @rdlaing: My take:Clinton: Let me explain about the emails   Press: Liar liar liar   Trump: I lie, its what I do.   Press: Ok"
CailleachSila|ericgarland|0.6908|0.0|0.769|0.231|"RT @ericgarland: IF on the off chance, Trump actually (and who could guess this) wins, then...wow, they've got quite an opening."
meghanchel|kurteichenwald|0.126|0.146|0.687|0.167|"RT @kurteichenwald: Putin staff consultant re: Trump choices: ""This is a fantastic team!""Remember when Romney said Russia biggest threat?"
daxis_gaming|RamonaCallender|0.4019|0.0|0.903|0.097|@RamonaCallender and yes it isn't that date yet so trump might not be the potus if you now abit more than the average person about elections
TCoop6231|deweydiva1|-0.1027|0.155|0.708|0.137|@deweydiva1 @MattMackowiak The specific claim I heard was that Trump is bad because he skips some intelligence brie https://t.co/diQkAErD4O
TCoop6231|twitter|-0.1027|0.155|0.708|0.137|@deweydiva1 @MattMackowiak The specific claim I heard was that Trump is bad because he skips some intelligence brie https://t.co/diQkAErD4O
cheapskare|goldengateblond|0.3818|0.0|0.88|0.12|RT @goldengateblond: Donald Trump's last press conference was July 27. He said he hoped Russia could find Hillary's emails. https://t.co/r4
cheapskare|t|0.3818|0.0|0.88|0.12|RT @goldengateblond: Donald Trump's last press conference was July 27. He said he hoped Russia could find Hillary's emails. https://t.co/r4
NickKilstein|BrendanNyhan|-0.4588|0.148|0.852|0.0|"RT @BrendanNyhan: At some point, Trump admin will act on this kind of rhetoric. Our democracy is in serious trouble if patriots do not spea"
born2fly2009|youtube|-0.7865|0.409|0.591|0.0|CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia https://t.co/pPQyxcSolP
RAOCES|tlaustin|-0.8074|0.316|0.684|0.0|"RT @tlaustin: @Hardees @Budweiser Your CEO as Trump's Sec of Labor is a disgusting offense against human decency. Puzder hates workers, wan"
nancy73gg|LindaSuhler|0.0|0.0|1.0|0.0|"RT @LindaSuhler: With PEOTUS Donald Trump we are reminded of when our Nation made these choices over 50 yrs ago, in Reagan's ""A Time For Ch"
MyGillianWill|mtaibbi|0.0|0.0|1.0|0.0|RT @mtaibbi: Fact: Donald Trump blasted both Ted Cruz and Hillary Clinton for their ties to Goldman. And he now has three Goldman vets in k
tibbidoe|SeabreezeCheryl|-0.2808|0.172|0.71|0.118|"RT @SeabreezeCheryl: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/ufmcVURB1v via @Bipart"
tibbidoe|bipartisanreport|-0.2808|0.172|0.71|0.118|"RT @SeabreezeCheryl: BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/ufmcVURB1v via @Bipart"
reroll|tfgnews)And|-0.6908|0.275|0.725|0.0|Retweeted Trump News Global (@tfgnews):And the execution should happen within 1 week of the crime. No more... https://t.co/C3E7BgfpVV
reroll|facebook|-0.6908|0.275|0.725|0.0|Retweeted Trump News Global (@tfgnews):And the execution should happen within 1 week of the crime. No more... https://t.co/C3E7BgfpVV
gant1014|Bipartisan|-0.2808|0.18|0.695|0.124|"BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/pJ2y2vUpSR via @Bipartisan Report"
gant1014|bipartisanreport|-0.2808|0.18|0.695|0.124|"BREAKING: Donald Trump Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) https://t.co/pJ2y2vUpSR via @Bipartisan Report"
neptune7321|floridaguy267|0.0|0.0|1.0|0.0|RT @floridaguy267: COAL Country Voting: Elliot County KY.  Registration 85% Democrat 8% GOP.  TRUMP 73% Hillary 27%.
Pikatyr|npfandos|0.2023|0.0|0.909|0.091|RT @npfandos: McCain urging a bipartisan reaction to hacking reports: You cant make this issue partisan. Its too important https://t.c
Pikatyr||0.2023|0.0|0.909|0.091|RT @npfandos: McCain urging a bipartisan reaction to hacking reports: You cant make this issue partisan. Its too important https://t.c
grandpooba5440|ianbremmer|-0.7089|0.237|0.763|0.0|RT @ianbremmer: Trump ignoring CIA evidence on Russian hacking for political expedience is the most irresponsible decision he has taken to
quebryant|trump_woman|-0.296|0.109|0.891|0.0|"RT @trump_woman: Report: Obama Wants to Become UN Secretary General, Netanyahu Doing Everything He Can to Stop Him https://t.co/toLjrt3Mdp"
quebryant|townhall|-0.296|0.109|0.891|0.0|"RT @trump_woman: Report: Obama Wants to Become UN Secretary General, Netanyahu Doing Everything He Can to Stop Him https://t.co/toLjrt3Mdp"
LaVerneWright13|AdamsFlaFan|-0.3612|0.167|0.739|0.094|"RT @AdamsFlaFan: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/wokIcX3tph via @crooksandliars"
LaVerneWright13|crooksandliars|-0.3612|0.167|0.739|0.094|"RT @AdamsFlaFan: Trump Okay With Pay-To-Play For Himself, Not Hillary Clinton | Crooks and Liars https://t.co/wokIcX3tph via @crooksandliars"
jennifer4nm|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
Sharonscofield2|WillBlackWriter|0.3182|0.0|0.897|0.103|RT @WillBlackWriter: Please tweet and ask your followers to tweet this Vine of Donald Trump asking Russia to hack Clinton. #Treasonhttps
pultuskpa|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
pultuskpa|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
AdamHeatherly|ChristophSouza|0.4728|0.126|0.627|0.247|@ChristophSouza @VitruvianMonkey oh yeah he was almost as bad with twitter as donald trump again midnights edge great videos
tomkardon|thehill|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
tomkardon|twitter|-0.8271|0.442|0.558|0.0|RT @thehill: Reporter who broke Watergate story calls Trump's lies worse than Nixon'shttps://t.co/LO4hyPAgxo https://t.co/mjJvsj5okk
TC_Stark|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
johnyc46|twitter|0.4215|0.0|0.843|0.157|Trump as a non politician did something McCain never could or will accomplish. Got Elected President. https://t.co/zLYOJk3VnS
HilaryVervers|bornmiserable|-0.1531|0.127|0.773|0.1|"RT @bornmiserable: Donald Trump, who literally begged Russia to find Hillary Clinton's emails, denies Russia's involvement in helping him w"
defendfreespeak|hawaiianlove68|0.7478|0.0|0.783|0.217|RT @hawaiianlove68: OMG what's it going to take to protect us from Trump and his minions? If anyone can say they aren't TERRIFIED RIGHT NOW
RachelK1967|AlwaysThinkHow|0.4767|0.0|0.853|0.147|RT @AlwaysThinkHow: #HolyShit Kellyanne Conway says Trump is going to put his own people in the intelligence community https://t.co/v3xjp
RachelK1967|t|0.4767|0.0|0.853|0.147|RT @AlwaysThinkHow: #HolyShit Kellyanne Conway says Trump is going to put his own people in the intelligence community https://t.co/v3xjp
mintyayaan|JoshButler|0.0|0.0|1.0|0.0|"RT @JoshButler: The New York Times piece on Australia's refugee policy is blistering. Dutton is our ""little Trump""  https://t.co/hvwnJ7XV7O"
mintyayaan|mobile|0.0|0.0|1.0|0.0|"RT @JoshButler: The New York Times piece on Australia's refugee policy is blistering. Dutton is our ""little Trump""  https://t.co/hvwnJ7XV7O"
JeremiahHope29|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
heliotactic|pdbuckland|0.4019|0.0|0.863|0.137|RT @pdbuckland: Yes. Actually they do. A lot of them. A HUUUUGE percentage of scientists. The @merchantsdoubt know it too.https://t.co/dLi
Mandari25733571|matthewjdowd|0.0|0.0|1.0|0.0|"RT @matthewjdowd: So Trump knows more about business than Wall Street Journal, more about military than Generals, and more about intelligen"
ValerieEllenLe1|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: Ltr from Hon Elijah Cummings asking Chaffetz to Investigate Trump biz conflicts#cnn #msnbc #AMJoy #cnnsotu #this
therightsarah|ElliottRHams|-0.1779|0.075|0.925|0.0|RT @ElliottRHams: .@Evan_McMullin has gone off the rails. Accusing Trump of disloyalty to America is too far even with the facts accounted
Jamiebalbier|davidfrum|0.2263|0.0|0.913|0.087|"RT @davidfrum: Its true that Donald Trump doesnt have a lot of foreign policy experience, but at least hes surrounded by knowledgeable p"
w_96_anthony|_joshjones1993|0.4404|0.0|0.408|0.592|@_joshjones1993 easy trump.
Fredio|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
scoutinfinity|Jodzio|-0.8625|0.346|0.654|0.0|"RT @Jodzio: Putin must have 'smoking gun"" that can ruin Trump. Probably sex related. But worse than anything that has been exposed so far."
IandPangurBan|aravosis|-0.6395|0.25|0.642|0.107|"RT @aravosis: And mind you, anonymous sources were more than good enough for Trump's racist conspiracy theories. But CIA sources on Russia?"
chefdnel|StopPC101|-0.34|0.224|0.658|0.118|@StopPC101 @realDonaldTrump Trump is an embarrassment who only ran to stoke his ego has no desire to govern
theshoewife|thedailybeast|0.0|0.0|1.0|0.0|"RT @thedailybeast: ""Hidden Figures"" is the movie Trump's America needs to see:  https://t.co/zBuYf87p2I https://t.co/R4qz0wQWha"
theshoewife|thedailybeast|0.0|0.0|1.0|0.0|"RT @thedailybeast: ""Hidden Figures"" is the movie Trump's America needs to see:  https://t.co/zBuYf87p2I https://t.co/R4qz0wQWha"
TAFORU|leahmcelrath|-0.3412|0.112|0.888|0.0|RT @leahmcelrath: NYTimes Editorial Board takes a stand &amp; even calls Trump out for not supporting an investigation into Russia hackinghttp
hgreenberg1|TeaPainUSA|0.0516|0.086|0.822|0.092|RT @TeaPainUSA: Is there any doubt left as to why Donald Trump won't release his tax returns?  Red Don needs to come clean or concede.  #Tr
ForestKing5280|theguardian|0.5859|0.0|0.798|0.202|Rex Tillerson: an appointment that would confirm Putin's US election win | US news | The Guardian https://t.co/qRxjiuQa1X
gaydaysLA|JuddLegum|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
gaydaysLA|medium|0.2023|0.0|0.917|0.083|"RT @JuddLegum: 1. John Bolton, according to Trump, has been one of his top foreign policy advisers from the outset https://t.co/oRUPSkz7NV"
Drewberedo|mateagold|-0.296|0.121|0.879|0.0|RT @mateagold: No president in recent history has filled a Cabinet with so many major donors. https://t.co/BbnJC608JZ https://t.co/zX9UKLSL
Drewberedo|washingtonpost|-0.296|0.121|0.879|0.0|RT @mateagold: No president in recent history has filled a Cabinet with so many major donors. https://t.co/BbnJC608JZ https://t.co/zX9UKLSL
LilleyDennese|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
LilleyDennese||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
vidaligodude|MartinWiener|-0.4767|0.147|0.853|0.0|@MartinWiener @AnthonyEinzig @realDonaldTrump prove me wrong. What would you call his business meetings abroad? All Trump biz thru POTUS.
wonderfullone|browntom1234|-0.4404|0.162|0.838|0.0|RT @browntom1234: @wonderfullone I imagine Alts are furiously making Joe-in-the-gas-chamber Pepe-Trump memes in Moms' basements the whole w
Sailfish157|BlackBelted|-0.7089|0.269|0.731|0.0|RT @BlackBelted: NBC having a fiduciary relationship with the president is completely unacceptable. Tell them to Dump Trump:  https://t.co/
Sailfish157|t|-0.7089|0.269|0.731|0.0|RT @BlackBelted: NBC having a fiduciary relationship with the president is completely unacceptable. Tell them to Dump Trump:  https://t.co/
mowser1970|FoxNews|0.5423|0.0|0.774|0.226|RT @FoxNews: Trump: We're Going to Start Saying 'Merry Christmas' Again https://t.co/rFmwtKQXIZ https://t.co/PexEqzNo9E
mowser1970|insider|0.5423|0.0|0.774|0.226|RT @FoxNews: Trump: We're Going to Start Saying 'Merry Christmas' Again https://t.co/rFmwtKQXIZ https://t.co/PexEqzNo9E
ArtOfSamWood|mattdpearce|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
ArtOfSamWood|mobile|0.0|0.0|1.0|0.0|"RT @mattdpearce: Behold, the next four years of our lives: https://t.co/fxANTMHByO https://t.co/oDbqsZLMOX"
Franco_AaronR|SenSanders|0.4767|0.08|0.691|0.229|"RT @SenSanders: I challenge Mr. Trump to tell the American people he'll keep his promises and veto cuts to Social Security, Medicare and Me"
jjen64|ClydeHaberman|-0.296|0.091|0.909|0.0|"RT @ClydeHaberman: Trump team says he had 1 of ""biggest Electoral College victories in history."" In fact, his % of electors puts him No. 46"
TheRealSusanA1|madworldnews|-0.6908|0.363|0.637|0.0|"NY Muslim Claims 3 White 'Trump' Fans Attacked Her, There's 1 Big Problem https://t.co/K9jMrZQVYA"
wakeupworldblog|change|0.8633|0.0|0.652|0.348|IT'S VERY IMPORTANT FOR THE AMERICAN PEOPLE TO KNOW FOR SURE THAT THE NEXT POTUS HAS BEEN ELECTED FAIR AND... https://t.co/kDw7bbDcko
DeborahWinchell|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
DaveJRosas|mikandynothem|-0.5267|0.167|0.833|0.0|RT @mikandynothem: President-elect Trump and our Police Officers will be working together again after a sickening Anti-Cop President.   #Bl
Deemoney521|JulieAnnLily|-0.3818|0.106|0.894|0.0|RT @JulieAnnLily: @robreiner We need emergency filing to halt EC. We have Russia interference &amp; collusion w trump &amp; trump team and GOP lead
moskaezul|DENVERSMKC|0.0|0.0|1.0|0.0|"RT @DENVERSMKC: Trump Inc makes $14.6M off of Trump running for President,how convenient and how unprecedented.I thought he was going to cl"
Ptmurf1016|FrankLuntz|0.0|0.0|1.0|0.0|"RT @FrankLuntz: ""How do you brief a president who refuses to believe what you tell him?""https://t.co/W2vLESP6l2"
Ptmurf1016|politico|0.0|0.0|1.0|0.0|"RT @FrankLuntz: ""How do you brief a president who refuses to believe what you tell him?""https://t.co/W2vLESP6l2"
YourAnonCentral|DrHaque|0.0|0.0|1.0|0.0|Democracy doesn't trump human rights. @DrHaque
17ninetyone|MattOrtega|0.0|0.0|1.0|0.0|RT @MattOrtega: Trump does it and *crickets* from the Republican leadership.Paul Ryan released a statement within nanoseconds after the C
princesseakitty|Womanista|0.5574|0.0|0.806|0.194|RT @Womanista: 'Teen Vogue' Writer @LaurenDuca Receives National Praise for Piece on Donald Trump https://t.co/HdR8x82h8Y https://t.co/9Ufs
princesseakitty|womanista|0.5574|0.0|0.806|0.194|RT @Womanista: 'Teen Vogue' Writer @LaurenDuca Receives National Praise for Piece on Donald Trump https://t.co/HdR8x82h8Y https://t.co/9Ufs
katieissweet_99|Tnacity|0.6145|0.0|0.851|0.149|@Tnacity @Al_Gorelioni @CNN Havent seen BS from Trump yet. Will b the 1st 2 say so if I did. And YES! People who know how 2 make money!#MAGA
mccurriel|OhEmmeG|0.128|0.0|0.87|0.13|RT @OhEmmeG: BREAKING: Trump announces Mojo Jojo as Secretary of Defense
sorenmacbeth|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
sorenmacbeth||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
charlesmire|afreedma|0.1531|0.0|0.89|0.11|"RT @afreedma: Trump falsely claims that ""nobody knows"" if global warming is real https://t.co/RcgsNAPCPf"
charlesmire|mashable|0.1531|0.0|0.89|0.11|"RT @afreedma: Trump falsely claims that ""nobody knows"" if global warming is real https://t.co/RcgsNAPCPf"
serge_poznanski|bloomberg|-0.34|0.179|0.821|0.0|business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/IkLASsHHyS https://t.co/KDKPsZJrcG
actionpollock|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
ChaosApathy|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
ChaosApathy|thegatewaypundit|0.0|0.0|1.0|0.0|RT @JackPosobiec: FBI Investigates Cybercrimes Not CIA I Told You That https://t.co/EThVy7qy45
Tamaraciocci|DavidCornDC|-0.7634|0.252|0.703|0.045|RT @DavidCornDC: Donald Trump appointing John Bolton shows that Trump was not serious in his post-invasion criticism of the Iraq war: https
ActionTime|ActionTime|0.8455|0.0|0.663|0.337|RT @ActionTime: Please Retweet:All US Security Agencies Should FULLY Brief Every Member of Electoral College on How Russia Helped Trump WON
WhoIsKeahJai|alwaystheself|0.0|0.0|1.0|0.0|RT @alwaystheself: Black folks at the beginning of 2016. Black folks at the end of 2016.Because black don't crack -- not even for Donal
DonMcKenzie|Delo_Taylor|-0.4019|0.124|0.876|0.0|RT @Delo_Taylor: Wikileaks is not the only spot for document dumps. Apparently nobody had the goods on Trump.  @mypostdemise @commietantric
C_BOYCE|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
C_BOYCE|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
cgbeige|ericgarland|-0.2052|0.114|0.805|0.08|"RT @ericgarland: And now, it's December 11th. Trump says he don't need no stinkin' intel agencies. Russia (BWA HAHAHAHAAAA) blames Ukrain"
KandiRider|porthos4424|0.296|0.0|0.855|0.145|"RT @porthos4424: Yeah, the Russians elected Donald Trump of President, on planet Hillary. https://t.co/NjqZXZ4jwW"
KandiRider|twitter|0.296|0.0|0.855|0.145|"RT @porthos4424: Yeah, the Russians elected Donald Trump of President, on planet Hillary. https://t.co/NjqZXZ4jwW"
clubfloozy|alwaystheself|0.0|0.0|1.0|0.0|RT @alwaystheself: Black folks at the beginning of 2016. Black folks at the end of 2016.Because black don't crack -- not even for Donal
beekuzz|JohnFugelsang|-0.2263|0.087|0.913|0.0|RT @JohnFugelsang: Trump blocks #millionwomanmarch from Lincoln Memorial despite the fact that the LM is actually owned by Americans who pa
MoMan60|sarahkendzior|-0.0258|0.196|0.613|0.19|RT @sarahkendzior: US Intelligence agencies fear reprisals over Russia revelations https://t.co/PP9qzrbB3s https://t.co/qwwUMIs3rV
MoMan60|theguardian|-0.0258|0.196|0.613|0.19|RT @sarahkendzior: US Intelligence agencies fear reprisals over Russia revelations https://t.co/PP9qzrbB3s https://t.co/qwwUMIs3rV
zoegits|washingtontimes|0.0|0.169|0.663|0.169|"Donald Trump-Tsai Ing-wen phone call raises hopes, fears in Taiwan - Washington Times https://t.co/4XFrMiZKUq"
Tstephenson23|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
Tstephenson23|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
thunderstruckcp|Tea4gunsSC|0.358|0.118|0.699|0.183|"@Tea4gunsSC Nobody did nothing til Trump, is that it? LOL! So, what's Trump's plan 2 deal with the deficit?"
campbellrock|MichaelGaree|-0.5267|0.204|0.739|0.057|"RT @MichaelGaree: Something comrade Trump's inner circle might want to consider: If he's charged with treason, guess who becomes co-conspir"
Myshiloh|davebernstein|-0.2808|0.151|0.746|0.104|"RT @davebernstein: BREAKING: Donald Trump, Mitch McConnell and James Comey Hit With TREASON Filing Monday Morning, Get Ready (DETAILS) http"
reblredhed|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
DanielHuculak|SarcasticHoney|-0.7269|0.243|0.757|0.0|RT @SarcasticHoney: @UniteAlbertans I suspect he is trying to distance himself from the Trump comparison as it is frankly media death.   @P
Dimipace|markwellsrector|0.4215|0.0|0.851|0.149|RT @markwellsrector: In Oct. Trump promoted a story that was a Russian state-controlled media fabrication. After being briefed. https://t.
Dimipace||0.4215|0.0|0.851|0.149|RT @markwellsrector: In Oct. Trump promoted a story that was a Russian state-controlled media fabrication. After being briefed. https://t.
inf0rmationist|thehill|0.0|0.0|1.0|0.0|RT @thehill: Christie turned down several positions in Trump administration: reporthttps://t.co/Ff4dxZ0zkz https://t.co/LVefpPfmiC
inf0rmationist|twitter|0.0|0.0|1.0|0.0|RT @thehill: Christie turned down several positions in Trump administration: reporthttps://t.co/Ff4dxZ0zkz https://t.co/LVefpPfmiC
polithist|EstherYuHsiLee|0.0|0.0|1.0|0.0|Trump gloats over Blacks who did not turn out to vote by @EstherYuHsiLee https://t.co/Mwzeq2WwBW
polithist|medium|0.0|0.0|1.0|0.0|Trump gloats over Blacks who did not turn out to vote by @EstherYuHsiLee https://t.co/Mwzeq2WwBW
jigokumimi|NBCNews|0.7579|0.0|0.698|0.302|"RT @NBCNews: CIA concludes Russia mounted covert operation to help Trump win, congressional official says https://t.co/hHlhMGJgwL https://t"
jigokumimi|nbcnews|0.7579|0.0|0.698|0.302|"RT @NBCNews: CIA concludes Russia mounted covert operation to help Trump win, congressional official says https://t.co/hHlhMGJgwL https://t"
kitten_nc|Dominus_Veritas|-0.357|0.262|0.738|0.0|RT @Dominus_Veritas: Ain't that grand? #MAGA #TRUMP https://t.co/hBOWKugJme
kitten_nc|twitter|-0.357|0.262|0.738|0.0|RT @Dominus_Veritas: Ain't that grand? #MAGA #TRUMP https://t.co/hBOWKugJme
bdanaher17|Reuters|0.2732|0.0|0.84|0.16|Rick Perry a leading candidate for U.S. energy post: source https://t.co/p9ysFp0dZo via @Reuters
bdanaher17|linkis|0.2732|0.0|0.84|0.16|Rick Perry a leading candidate for U.S. energy post: source https://t.co/p9ysFp0dZo via @Reuters
Rickeyleetw|vivelafra|-0.5622|0.251|0.624|0.125|RT @vivelafra: THE RUSSIA HOAX: Julian Assange acknowledges murdered DNC staffer Seth Rich was Wikileaks' source.  Why is MSM covering this
ThelmaOAgyekum|CNN|0.0772|0.0|0.902|0.098|"RT @CNN: Trump on cabinet picks: ""I want people that made a fortune"" https://t.co/w9ZXsRxORA"
ThelmaOAgyekum|snappytv|0.0772|0.0|0.902|0.098|"RT @CNN: Trump on cabinet picks: ""I want people that made a fortune"" https://t.co/w9ZXsRxORA"
lanorte1|JohnCena|0.0|0.0|1.0|0.0|". @JohnCena looks at the world through @realDonaldTrumps eyes on ""SNL""  by @lee_moran https://t.co/hPajSH8jmg via @HuffPostComedy"
lanorte1|huffingtonpost|0.0|0.0|1.0|0.0|". @JohnCena looks at the world through @realDonaldTrumps eyes on ""SNL""  by @lee_moran https://t.co/hPajSH8jmg via @HuffPostComedy"
sherrilee7|MichaelGaree|-0.5267|0.204|0.739|0.057|"RT @MichaelGaree: Something comrade Trump's inner circle might want to consider: If he's charged with treason, guess who becomes co-conspir"
KarmaKittySays|vivelafra|-0.6486|0.194|0.806|0.0|"RT @vivelafra: BIG 6: After criminally colluding with his opponent for 18 months, MSM is now trying to suggest #Trump had an unfair advanta"
princessmom122|KaylinWinters2|-0.8271|0.386|0.614|0.0|RT @KaylinWinters2: GOP was willing to prosecute Hillary Clinton for fake scandals &amp; lies but evidence of trump colluding with Russia? Not
DangerVenture|newyorker|0.6705|0.0|0.353|0.647|The best closing sentence. https://t.co/LhAfu9yo5o
jimi_jimijones|ANDtwenty1|0.765|0.0|0.515|0.485|@ANDtwenty1 if trump can win he def can lol
RandallBeard88|Cernovich|0.103|0.079|0.787|0.134|"RT @Cernovich: Trump is not a perfect man, flawed to be sure like everyone else, but compared to Clintons (either of them), he's a saint."
starfishncoffee|goldengateblond|0.9423|0.0|0.435|0.565|"RT @goldengateblond: Easy to laugh at Trump's ""I'm, like, smart"" comment, but claiming divine intelligence isn't just narcissistic. That's"
mariean24614777|YouTube|0.0772|0.161|0.657|0.182|President-Elect Trump Is Tweeting To Relieve The Pressure https://t.co/FbM4dO73WF via @YouTube
mariean24614777|youtube|0.0772|0.161|0.657|0.182|President-Elect Trump Is Tweeting To Relieve The Pressure https://t.co/FbM4dO73WF via @YouTube
gayginsburned|softbutchkate|0.6633|0.0|0.67|0.33|"RT @softbutchkate: YEAHHHH ALEC WON FOR TRUMP, TAKE THAT @realDonaldTrump"
cocktailgurl17|Khanoisseur|-0.4588|0.15|0.85|0.0|RT @Khanoisseur: 2 reasons for trump rejecting daily intel briefings:1. Plausible deniability2. Busy making side deal$$ for himself @mrp
ActionTime|ActionTime|0.3182|0.0|0.892|0.108|RT @ActionTime: Please Retweet: Presidential Ethics Counsel: How Can Trump Regulate Financial Sector When He Owes Millions To Banks? https:
penguingotico|jeongshk|-0.296|0.167|0.833|0.0|RT @jeongshk: No bangtao temostemertrumpduas dilmas lulaTo sentindo q isso est politicamente errado
killjoykittens1|RalfThePowerful|-0.2023|0.083|0.917|0.0|"RT @RalfThePowerful: When confronted with evidence that Russia worked to elect him, rather than ""I can't be bought,"" Trump's statement was"
pennylane314|ELCALBO1961|0.0|0.0|1.0|0.0|@ELCALBO1961 @KellyannePolls how much you wanna bet she is fuckin trump
IntrepidCommute|on2_off4|0.4836|0.184|0.668|0.148|"RT @on2_off4: obama doesn't want Trump ""whining""...I guess it cuts into what barry does best and he doesn't want competition! ""bush did it!"
BuffyMaxSFCA|aravosis|-0.765|0.355|0.645|0.0|"RT @aravosis: I still cant decide if Trump is a liar, an idiot, or delusional. https://t.co/Z2VlmbuRf8"
BuffyMaxSFCA|twitter|-0.765|0.355|0.645|0.0|"RT @aravosis: I still cant decide if Trump is a liar, an idiot, or delusional. https://t.co/Z2VlmbuRf8"
Redrebel92|twitter|0.0|0.0|1.0|0.0|Release your tax returns Mr. Trump!!!! https://t.co/cqEIxfmREW
Nazaninstyle|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Nazaninstyle||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
jaystebbins|sluggahjells|-0.5216|0.128|0.872|0.0|"RT @sluggahjells: In which Trump comes to the Army-Navy game, only to then diss the Army-Navy game about not having the ""best football."" ht"
grandpooba5440|RVAwonk|-0.3818|0.185|0.725|0.091|RT @RVAwonk: Bottom line: The FBI and CIA agree that Russia hacked our democratic process. So why is #Trump still denying Russian interfere
AfricaOhAfrica2|stanleyrogouski|-0.1027|0.174|0.714|0.112|RT @stanleyrogouski: Do the Democrats actually believe they're going to stop Trump by accusing him of being a Russian asset?
abelmezg|canalN_|-0.296|0.18|0.82|0.0|"@canalN_ seor Trump, no olvides que America es para los Americanos."
4joycie|npfandos|0.4515|0.0|0.835|0.165|"@npfandos does this trump person have a crystal ball?  is he capable of ""knowing things"" by osmosis?"
KPMcClave|DanRather|0.3612|0.0|0.894|0.106|RT @DanRather: Actually people do know climate change is real - like scientists and almost every other head of state in the world.https:/
SNUGSFBay|adambosworth|-0.5267|0.298|0.702|0.0|RT @adambosworth: Trumps Threat to the Constitution - https://t.co/U6QpjsgsYB https://t.co/643AAm9OO4
SNUGSFBay|nytimes|-0.5267|0.298|0.702|0.0|RT @adambosworth: Trumps Threat to the Constitution - https://t.co/U6QpjsgsYB https://t.co/643AAm9OO4
MissUSA56|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
MissUSA56|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
haarusso|au48|-0.2263|0.192|0.808|0.0|Trump hints he's still undecided about Tillerson | #RexTillerson https://t.co/nImBHGqDfJ
debinny55|AdamSmith_usa|0.0|0.0|1.0|0.0|RT @AdamSmith_usa: This fleece has more experience than Donald Trump. https://t.co/USGojcf5lX
debinny55|twitter|0.0|0.0|1.0|0.0|RT @AdamSmith_usa: This fleece has more experience than Donald Trump. https://t.co/USGojcf5lX
jaggy123|McClatchyDC|0.5859|0.0|0.826|0.174|"RT @McClatchyDC: Since his election win, Trump has talked to Putin more than any other world leader https://t.co/mLBJ0589N3 https://t.co/QN"
jaggy123|mcclatchydc|0.5859|0.0|0.826|0.174|"RT @McClatchyDC: Since his election win, Trump has talked to Putin more than any other world leader https://t.co/mLBJ0589N3 https://t.co/QN"
Mary8941|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
serenityatsea|funder|0.0|0.0|1.0|0.0|"RT @funder: #TRUMPLEAKS Donald &amp; Ivanka Trump sent 1,347 shipments for clothing line w/Iranian affiliated cos #GrabYourWallet #amjoy @JoyAn"
damienics|Noahpinion|-0.6124|0.263|0.647|0.091|"RT @Noahpinion: Prediction: Trump will push hard to kill alternative energy technology. After all, Russia is a petrostate... https://t.co/f"
damienics|twitter|-0.6124|0.263|0.647|0.091|"RT @Noahpinion: Prediction: Trump will push hard to kill alternative energy technology. After all, Russia is a petrostate... https://t.co/f"
goddesslaney|TheDailyEdge|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
goddesslaney|twitter|-0.3612|0.181|0.7|0.119|RT @TheDailyEdge: I think Paul Ryan's enthusiasm for killing Medicare may be blinding him to some of Trump's flaws. https://t.co/ZfCi71ykKN
SharonS72105601|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
SharonS72105601|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
pol_quebec|lapresse|-0.4939|0.176|0.824|0.0|Trump menace de ne plus reconnatre le principe de la Chine unique https://t.co/zHGvSpchIe #polqc #assnat https://t.co/OUtddjWvZ3
bighungrygeek|JoyAnnReid|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
bighungrygeek|twitter|0.3818|0.0|0.794|0.206|"RT @JoyAnnReid: A unified theory of Trump, Putin and Exxon Mobil. https://t.co/tLUFgAep9r"
HonkyTonkNights|breitbart|0.4939|0.0|0.758|0.242|Five Actions President Trump Can Take to Save 2nd Amendment https://t.co/p9T67ynOAM
Mc_Heckin_Duff|ericgarland|-0.2052|0.114|0.805|0.08|"RT @ericgarland: And now, it's December 11th. Trump says he don't need no stinkin' intel agencies. Russia (BWA HAHAHAHAAAA) blames Ukrain"
ProgressiveJill|MayorHodges|0.529|0.0|0.784|0.216|"RT @MayorHodges: Today I joined @ChicagosMayor in urging President-elect Trump not to cut DACA, which helps immigrant children. https://t.c"
ProgressiveJill||0.529|0.0|0.784|0.216|"RT @MayorHodges: Today I joined @ChicagosMayor in urging President-elect Trump not to cut DACA, which helps immigrant children. https://t.c"
granbulls|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
granbulls|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
wildwonderweb|sarahkendzior|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
wildwonderweb|twitter|0.1027|0.115|0.752|0.133|RT @sarahkendzior: Elizabeth Warren is calling for an audit of Trump's finances due to conflicts of interest #Resist https://t.co/HPS5Xiank9
triplesss1001|tomtomorrow|-0.3182|0.182|0.704|0.114|"RT @tomtomorrow: Trump's  victory is as if your loved one died, and you grieve, and then they are brought back to life the next day and kil"
macmcd|starfirst|-0.6908|0.305|0.695|0.0|RT @starfirst: @deejay90192 Donald Trump and the Republican's leaders are guilty of treason. They're  traitors
AvaSimon1984|TheDailyShow|0.0772|0.118|0.749|0.134|RT @TheDailyShow: .@jordanklepper checks out the first stop on Donald Trumps Thank You Tour. https://t.co/RCcCU3dZb7 https://t.co/DXHCRP
AvaSimon1984|cc|0.0772|0.118|0.749|0.134|RT @TheDailyShow: .@jordanklepper checks out the first stop on Donald Trumps Thank You Tour. https://t.co/RCcCU3dZb7 https://t.co/DXHCRP
Fire_Badger|CoolCalmCam|0.1774|0.108|0.751|0.141|@CoolCalmCam holy shit r/politics is nothing but shitting on trumpthis would get a lot of people hateswarmed 2 months ago
CaroleMyers|FBI=only|-0.2411|0.089|0.911|0.0|"Does beg the question, was Comey in cahoots wi/Russia to elect Trump? @FBI=only agency not sure R;s goal was electi https://t.co/hTS1r7nwU9"
CaroleMyers|twitter|-0.2411|0.089|0.911|0.0|"Does beg the question, was Comey in cahoots wi/Russia to elect Trump? @FBI=only agency not sure R;s goal was electi https://t.co/hTS1r7nwU9"
BerkowitzAnne|linkis|0.3818|0.0|0.729|0.271|Schwarzenegger Defends Trump's 'Celebrity Apprentice' Producer Credit https://t.co/PrGN0gqMaO
lnfoComunio|elpais|0.0|0.0|1.0|0.0|Va traicionar Trump a los trabajadores? https://t.co/Mnifgy2VTQ
BollmerJason|GrrrGraphics|0.0|0.0|1.0|0.0|RT @GrrrGraphics: New #BenGarrison #Cartoon #NewBroom #Trump #Maga Sweep away the dirt/ #FakeNews ! more cartoons at https://t.co/Oj98iIxEA
BollmerJason|t|0.0|0.0|1.0|0.0|RT @GrrrGraphics: New #BenGarrison #Cartoon #NewBroom #Trump #Maga Sweep away the dirt/ #FakeNews ! more cartoons at https://t.co/Oj98iIxEA
JJohnson2u|ProtestDaily|-0.2263|0.119|0.881|0.0|RT @ProtestDaily: #Protest #Trump Protesters decry President-Elect Trump on International Human Rights Day - KMSP-TV https://t.co/EwOjzovZ9E
JJohnson2u|fox9|-0.2263|0.119|0.881|0.0|RT @ProtestDaily: #Protest #Trump Protesters decry President-Elect Trump on International Human Rights Day - KMSP-TV https://t.co/EwOjzovZ9E
anthonyzenkus|Delo_Taylor|-0.3818|0.094|0.906|0.0|"RT @Delo_Taylor: If the goal was to keep Trump from ever becoming POTUS, the first thing you shoulda done was fight to keep HRC from being"
trulyguide|goldengateblond|0.4201|0.0|0.872|0.128|RT @goldengateblond: Absolutely agree. Speaking of other countries: Can we get your thoughts on the Trump/Putin situation? Haven't seen you
mowser1970|DaysOfTrump|-0.4215|0.132|0.818|0.05|RT @DaysOfTrump: .@SpeakerRyan We know #FakeNews &amp; #Russia hysteria are globalist attempt to prevent Trump from rebuilding our country. The
moralesdc|bmangh|0.6249|0.0|0.733|0.267|"RT @bmangh: Gen. Barry McCaffrey withdraws support of Trump national security advisor, calls for investigation https://t.co/RIJztQRROe"
moralesdc|m|0.6249|0.0|0.733|0.267|"RT @bmangh: Gen. Barry McCaffrey withdraws support of Trump national security advisor, calls for investigation https://t.co/RIJztQRROe"
eph4_15|washingtonpost|-0.4019|0.144|0.856|0.0|"Small SAMPLING of The Myriad of Conflicting Ideas coming from Donald ""Anti-Establishment"" Trump [Sarc] https://t.co/3KTkxYCh6G #PJNET #CCOT"
drandreaj|rudepundit|-0.765|0.248|0.752|0.0|"RT @rudepundit: Maybe Trump is too dumb to understand that the word ""intelligence"" isn't meant as an insult to those being briefed."
Brooke888888|Bros4Hillary|0.4404|0.0|0.633|0.367|RT @Bros4Hillary: Good for her.  https://t.co/Idm9vtGoXW
Brooke888888|buzzfeed|0.4404|0.0|0.633|0.367|RT @Bros4Hillary: Good for her.  https://t.co/Idm9vtGoXW
KatCeccotti|funder|0.8176|0.0|0.706|0.294|"RT @funder: Breaking: Ku Klux Klan parades in Roxboro, NC celebrating Trump win #cnn #msnbc #ncpol #amjoy #antitrump #trumpleaks https://t."
KatCeccotti||0.8176|0.0|0.706|0.294|"RT @funder: Breaking: Ku Klux Klan parades in Roxboro, NC celebrating Trump win #cnn #msnbc #ncpol #amjoy #antitrump #trumpleaks https://t."
milkyyoon_|jiyongal|-0.6841|0.188|0.812|0.0|RT @jiyongal: SEUNGHYUN MAKING HIS DISGUST FOR DONALD TRUMP KNOWN WITHOUT EVEN SAYING ANYTHING AT ALL IM SVRSMSIGNG WOKE KING https://t.co/
milkyyoon_|t|-0.6841|0.188|0.812|0.0|RT @jiyongal: SEUNGHYUN MAKING HIS DISGUST FOR DONALD TRUMP KNOWN WITHOUT EVEN SAYING ANYTHING AT ALL IM SVRSMSIGNG WOKE KING https://t.co/
Powder08|kurteichenwald|-0.5423|0.176|0.824|0.0|"RT @kurteichenwald: Fox/Cheney went nuts when found out Obama got intel briefings in writing, rather than read to him. But Trump no briefin"
FALSEKXNGG|CloudN9neSyrup|-0.7184|0.318|0.682|0.0|"RT @CloudN9neSyrup: She's talking nonsense but forget Trump and Hillary, this man Gary Johnson has no chill  https://t.co/DrJB0tvJda"
FALSEKXNGG|twitter|-0.7184|0.318|0.682|0.0|"RT @CloudN9neSyrup: She's talking nonsense but forget Trump and Hillary, this man Gary Johnson has no chill  https://t.co/DrJB0tvJda"
Newyorker2212|peglepetit|0.8445|0.062|0.582|0.356|RT @peglepetit: @KellyannePolls @nypost  churlish comment.  So hard for the winner to be gracious? Get Trump to #reimburseNYC for security
Bjb58barb|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Bjb58barb||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
mdufay|marklevinshow|-0.6369|0.276|0.724|0.0|RT @marklevinshow: More Goldman Sachs appointments; I thought Trump hated Goldman Sachs https://t.co/d93fhyI6cG
mdufay|conservativereview|-0.6369|0.276|0.724|0.0|RT @marklevinshow: More Goldman Sachs appointments; I thought Trump hated Goldman Sachs https://t.co/d93fhyI6cG
JBax52|MtnMD|0.34|0.0|0.888|0.112|RT @MtnMD: RT @JesseLehrich: a year ago today:  Trump's National Security Adviser sitting next to Putin at the @RT_com gala https://t.co/5q
JBax52|t|0.34|0.0|0.888|0.112|RT @MtnMD: RT @JesseLehrich: a year ago today:  Trump's National Security Adviser sitting next to Putin at the @RT_com gala https://t.co/5q
CarolJo76077222|Kosart20|-0.7885|0.351|0.552|0.098|RT @Kosart20: @thedailybeast you mean LYING. Trump keeps LYING about who is responsible for the hacking
ArgentinaPatito|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS:Memo:Ivanka Trump's Iranian shipments-all made while sanctions in place on Iran#GrabYourWallet #amjoy #msnbc #mon
dayadelreys|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
JennyMenezess|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
LDB3_Esquire|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
SheilaSmithCFR|fravel|0.0|0.0|1.0|0.0|"RT @fravel: ""Chinas senior foreign policy official, Yang Jiechi, met with Lt. Gen. Michael T. Flyn"" https://t.co/11OnQiEfAX"
SheilaSmithCFR|mobile|0.0|0.0|1.0|0.0|"RT @fravel: ""Chinas senior foreign policy official, Yang Jiechi, met with Lt. Gen. Michael T. Flyn"" https://t.co/11OnQiEfAX"
NancyLebMiller|LadyDoc4Trump|0.0|0.0|1.0|0.0|"RT @LadyDoc4Trump: Our ""president"" says NOTHING, NADA, ZERO about #Christian genocide by his Muslim brothers.#Trump speaks #Truth on it."
greatwallofsam|lauraolin|0.0|0.0|1.0|0.0|RT @lauraolin: Kirk Douglas turns 100 today. He was 16 when Hitler came to power. Here's what he thinks about Trump: https://t.co/DZ6PmDQux
greatwallofsam|t|0.0|0.0|1.0|0.0|RT @lauraolin: Kirk Douglas turns 100 today. He was 16 when Hitler came to power. Here's what he thinks about Trump: https://t.co/DZ6PmDQux
Tamaraciocci|JuddLegum|0.0|0.0|1.0|0.0|RT @JuddLegum: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/oRUPSkz7NV https:
Tamaraciocci|medium|0.0|0.0|1.0|0.0|RT @JuddLegum: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/oRUPSkz7NV https:
drcastillo55|WayneDupreeShow|-0.4767|0.171|0.829|0.0|RT @WayneDupreeShow: Rep. Tulsi Gabbard Says Democrats Wrong To Bash Trump For Retired General Picks https://t.co/62oDMIBBmO
drcastillo55|newsninja2012|-0.4767|0.171|0.829|0.0|RT @WayneDupreeShow: Rep. Tulsi Gabbard Says Democrats Wrong To Bash Trump For Retired General Picks https://t.co/62oDMIBBmO
SandraPitts14|funder|0.0|0.0|1.0|0.0|RT @funder: #TRUMPLEAKS: US Senators letter to Senate leaders-investigate Trump for Russian espionage#cnn #msnbc #AMJoy #cnnsotu #thiswee
katriord|ericgarland|0.5719|0.0|0.817|0.183|RT @ericgarland: Trump looks like he swallowed a goldfish and stares at the floor a bit too long.As if maybe a joke has gone too far.
Shirleyann27|misscherryjones|0.0|0.0|1.0|0.0|"RT @misscherryjones: Just when I think the CIA-Russia-Trump takes can't get any hotter, along comes John Bolton with a torch."
MissPride2u|USARedOrchestra|0.0|0.0|1.0|0.0|"RT @USARedOrchestra: CT Rep. Jim Himes call Trump ""completely unhinged"" and calls for the electoral college to do what it was designed for."
michaeljordaned|BCAppelbaum|0.0772|0.0|0.929|0.071|RT @BCAppelbaum: Trump most resembles the average American in the number of hours he spends watching television. https://t.co/4ynwJAWnzh
michaeljordaned|twitter|0.0772|0.0|0.929|0.071|RT @BCAppelbaum: Trump most resembles the average American in the number of hours he spends watching television. https://t.co/4ynwJAWnzh
MythicalStig|kurteichenwald|0.2263|0.087|0.791|0.123|"RT @kurteichenwald: Trump's approval rating now lower than all PRESIDENT averages except for 2nd term of Truman, Nixon and GW Bush. Unprece"
veevardhan|simonhelberg|0.8126|0.0|0.657|0.343|RT @simonhelberg: cool just go on instinct I'm sure there's not much to this whole president thing oh my god help https://t.co/uqnX4BatOq
veevardhan|medium|0.8126|0.0|0.657|0.343|RT @simonhelberg: cool just go on instinct I'm sure there's not much to this whole president thing oh my god help https://t.co/uqnX4BatOq
zenithguy|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
lyseee_|jdakwar|-0.8779|0.387|0.613|0.0|"RT @jdakwar: Horrific genocidal statement by military veteran and former congressman Allen West, a notorious Muslim hater emboldened by Tru"
ChiefG4LSU|RichardTBurnett|0.8316|0.0|0.63|0.37|RT @RichardTBurnett: Everything is coming back thanks to Donald Trump:1. Pride in America.2. Saluting American flag.3. Merry Christmas.
MiaShaw|washingtonpost|-0.4019|0.144|0.856|0.0|RT @washingtonpost: Trumps last press conference was where he asked Russia to release Clintons hacked emails https://t.co/epszMRvnDs
MiaShaw|washingtonpost|-0.4019|0.144|0.856|0.0|RT @washingtonpost: Trumps last press conference was where he asked Russia to release Clintons hacked emails https://t.co/epszMRvnDs
ValkyrieHanna7|JeannieM0625|0.0|0.0|1.0|0.0|@JeannieM0625 @AmericaNewsroom and p will get over it!  Thats normalizing Trump &amp; all of his disgustingness.  Theres nothing normal about it
cablefixer|danfelix82|0.0|0.0|1.0|0.0|@danfelix82  It's cause they weren't allowed to go to white schools.. Geez You're a total trump moron..
JP61926104|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
JP61926104|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
radiofreeorg|radiofree|0.0|0.0|1.0|0.0|Baltimore City Council members Defend Resolution Condemning Trump's Bigotry... https://t.co/vGmailQ3sS
rlswanson5|Run_IsHere|-0.5423|0.179|0.821|0.0|RT @Run_IsHere: Another Republican crook trying to cover up a crime against America by Russia and Trump. https://t.co/SPWm5dw1Gg
rlswanson5|twitter|-0.5423|0.179|0.821|0.0|RT @Run_IsHere: Another Republican crook trying to cover up a crime against America by Russia and Trump. https://t.co/SPWm5dw1Gg
jmpilon|MaggieJordanACN|0.5165|0.058|0.746|0.196|RT @MaggieJordanACN: Interesting point:Trump is not denying the hack.He's questioning WHO did the hack and WHO put out the story. https:
DMacOttawa|ezlusztig|-0.6249|0.17|0.83|0.0|"RT @ezlusztig: Purely on the basis of information publicly available - just the tip of an iceberg, presumably - Obama could devastate Trump"
zebedol|twitter|-0.5228|0.144|0.856|0.0|"And, of course, all the Republicans are yelling to impeach him.  When will this madness end? Go away, Trump.  Far a https://t.co/BWiVmFxXAf"
whitewolf8214|LouDobbs|-0.6597|0.221|0.779|0.0|RT @LouDobbs: The Ignorance of the Left is Rising to the Level of Sheer Madness #MAGA #Trump @FoxBusiness @FoxNews #Dobbs https://t.co/LTyu
whitewolf8214|t|-0.6597|0.221|0.779|0.0|RT @LouDobbs: The Ignorance of the Left is Rising to the Level of Sheer Madness #MAGA #Trump @FoxBusiness @FoxNews #Dobbs https://t.co/LTyu
sud_vijay|matthewjdowd|0.4019|0.0|0.886|0.114|"RT @matthewjdowd: Trump calling himself a ""smart person"" reminds me of margaret thatcher: ""if you have to tell people you are a lady, you p"
xBlade13710x|JoeySalads|0.5719|0.0|0.778|0.222|RT @JoeySalads: None of these Liberal celebs left the country yet after Trump won.
maddiecarey5187|sydneyhfluty|0.0|0.0|1.0|0.0|RT @sydneyhfluty: Maybe trump should build a wall between Mingo and Wayne 
karma1120|MelindaThinker|0.0|0.0|1.0|0.0|RT @MelindaThinker: Calls for a second election after Russia's meddling are increasing https://t.co/ESjr1JeEGl
karma1120|politicususa|0.0|0.0|1.0|0.0|RT @MelindaThinker: Calls for a second election after Russia's meddling are increasing https://t.co/ESjr1JeEGl
bbroom01|AngrySalmond|0.624|0.0|0.746|0.254|RT @AngrySalmond: 100 year-old Kirk Douglas takes down Donald Trump. Absolutely brilliant. https://t.co/rU5GGbDGwE
bbroom01|twitter|0.624|0.0|0.746|0.254|RT @AngrySalmond: 100 year-old Kirk Douglas takes down Donald Trump. Absolutely brilliant. https://t.co/rU5GGbDGwE
crime18458238|AJDelgado13|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
crime18458238|twitter|-0.0258|0.127|0.751|0.121|"RT @AJDelgado13: Well, what do we have here.... Put your pitchforks down, Trump critics. https://t.co/7BpFnPQGfD"
Tull007|saletan|0.4019|0.0|0.899|0.101|RT @saletan: Trump and aides went on TV to dismiss a CIA report they haven't seen. That's the story: They treat intel on Russian ops as a t
mimi_x4|laurine3215|0.5719|0.0|0.871|0.129|RT @laurine3215: Trump watches all news stations to see what they have to say about him. That's how he grades all media. He loves Fox and H
banreportcards|gmbutts|0.0|0.0|1.0|0.0|https://t.co/BbfePg05WH@gmbutts
banreportcards|medium|0.0|0.0|1.0|0.0|https://t.co/BbfePg05WH@gmbutts
andythibeault|RachaelRad|0.6808|0.145|0.597|0.258|RT @RachaelRad: The best smartest take I've read about this whole mess in awhile and it's out of the television critic section. https://t
andythibeault||0.6808|0.145|0.597|0.258|RT @RachaelRad: The best smartest take I've read about this whole mess in awhile and it's out of the television critic section. https://t
TimGOGOGomez|LOLGOP|-0.6917|0.248|0.67|0.082|RT @LOLGOP: Trump doesn't like to be known as the biggest popular vote loser to be elected in modern history. It would be rude to point tha
fraterrisus|Pinboard|-0.7783|0.281|0.719|0.0|"RT @Pinboard: Remember, if you work at Google or Facebook and frustrated by management inaction on Trump, leak to uncle Pinboard. 415 610 0"
JohnSil08042759|SenSanders|0.0|0.0|1.0|0.0|"RT @SenSanders: Mr. Trump may not know it, and his nominee for EPA administrator may not know it, but the debate is over. Climate change is"
ChristineAdams3|laureldavilacpa|0.0|0.0|1.0|0.0|RT @laureldavilacpa: #ImStillNotOver Before the election the Senate was briefed by the CIA of #RussianHackers electioneering for Trump - an
maropesa|NBCNews|0.0516|0.145|0.661|0.194|RT @NBCNews: A slap in the face. That's how intelligence agencies see Trump's rejection of findings on Russia https://t.co/k6QZxwjtem https
maropesa|nbcnews|0.0516|0.145|0.661|0.194|RT @NBCNews: A slap in the face. That's how intelligence agencies see Trump's rejection of findings on Russia https://t.co/k6QZxwjtem https
negilyn|EW|0.802|0.0|0.753|0.247|RT @EW: Do NOT tweet Donald Trump right now telling him that Alec Baldwin just won a #CriticsChoice award for his #SNL portrayal of him. 
pinklady404|DavidYankovich|-0.1531|0.158|0.739|0.102|RT @DavidYankovich: My immediate goal is stopping Trump.Then we are going to end the GOP for their treason of the US by supporting enemie
Mrsjagray|kurteichenwald|0.4215|0.0|0.887|0.113|"RT @kurteichenwald: Reminder of what I said in July, cause Ive known Trump since 87: Doesnt wanna BE prez, wants applause. Wont sit 4 brief"
WNHastings|AJUpFront|0.2023|0.129|0.679|0.193|"@AJUpFront @mehdirhasan Thanks for trying Mehdir.  Like you, we remember what Mr. Trump originally said and it was a total ban on Muslims."
JoshuaJrrp42|DavidBellCBC|0.0|0.0|1.0|0.0|@DavidBellCBC @Dfildebrandt Canada needs our own Daddy (Donald Trump)
mollylmaguire|AlwaysThinkHow|0.4767|0.0|0.853|0.147|RT @AlwaysThinkHow: #HolyShit Kellyanne Conway says Trump is going to put his own people in the intelligence community https://t.co/v3xjp
mollylmaguire|t|0.4767|0.0|0.853|0.147|RT @AlwaysThinkHow: #HolyShit Kellyanne Conway says Trump is going to put his own people in the intelligence community https://t.co/v3xjp
cxpey|AntTheIcon|0.4515|0.141|0.617|0.242|RT @AntTheIcon: worst 2 teams? 49ers with a BLM QB and the BROWNS. best record? the AMERICAN conference PATRIOTS whose QB publicly supports
SukiOshea|KellyannePolls|-0.296|0.121|0.879|0.0|@KellyannePolls @realDonaldTrump @andrewrcamp and Trump knows about public education ... How...? Must have missed that one. #notmypresident
menjicm|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
kbal3259|Diana25017037|-0.4003|0.233|0.614|0.153|RT @Diana25017037: @APPROVEMAN @LisaBloom @GloriaAllred @jillharth @thejessicadrake @danabrams  THANK YOU! NOBODY TALKS ABOUT THE VIOLENT T
Gjizzle55|AriMelber|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
Gjizzle55|t|-0.7717|0.355|0.645|0.0|"RT @AriMelber: Trump previously criticized Obama for missing intel briefings - inaccurate at the time, hypocritical now: https://t.co/301NA"
srauer20|blogdiva|0.3612|0.0|0.889|0.111|"RT @blogdiva: @brownblaze @leahmcelrath giuliani, like chris christie, was given the boot. they're guidos as far as Trump is concerned, and"
templvr|business|-0.34|0.167|0.833|0.0|RT @business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/6l8izhUs9D https://t.co/0drSTTUrnr
templvr|bloomberg|-0.34|0.167|0.833|0.0|RT @business: Japan watches uneasily as Trump shakes up Taiwan-China relations https://t.co/6l8izhUs9D https://t.co/0drSTTUrnr
venrala|TheDemocrats|0.0|0.0|1.0|0.0|"RT @TheDemocrats: ""When Trump said ""drain the swamp,"" he really just meant ""appoint a bunch of Goldman Sachs bankers."" https://t.co/8JnGFai"
venrala|t|0.0|0.0|1.0|0.0|"RT @TheDemocrats: ""When Trump said ""drain the swamp,"" he really just meant ""appoint a bunch of Goldman Sachs bankers."" https://t.co/8JnGFai"
FrankenFert|twitter|-0.8481|0.351|0.649|0.0|"Lmfaoooo that racist white man is shook over Trump and his recent actions. Bitch I'm dying, that nigga like........ https://t.co/LaVApmturc"
teraphin|StephenKing|-0.6249|0.227|0.773|0.0|RT @StephenKing: Trump's proposed cabinet is the worst in American history: a motley crew of plunder-monkeys.
Wyohawk|mitchellvii|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
Wyohawk|thegatewaypundit|0.128|0.123|0.726|0.151|RT @mitchellvii: FBI Investigation Refutes CIA=&gt; There's No Evidence Russia Tried to Help Trump https://t.co/Tvsa5cwA0W
anythingbutdem|twitter|0.4215|0.0|0.896|0.104|1) I'm a Republican. 2) I'm 32. 3) True. 4) We have yet to see if Trump is much of a Republican at all. All signs p https://t.co/IPCAY0hdhE
Newsstand_|nytimes|0.0|0.0|1.0|0.0|Trump Suggests Using Bedrock China Policy as Bargaining Chip - New York TimesNew York TimesTrump Suggests Usin https://t.co/rUCDPmHZEP
MikeMmwh|IngrahamAngle|0.5106|0.0|0.815|0.185|@IngrahamAngle Challenge for Trump: Facing a sea of lefty journalists and reporters who all think they are way smarter than he is...
TweeetBug|GoAngelo|0.2023|0.094|0.779|0.127|RT @GoAngelo: NBC has a financial stake in Trump's reputation. How can they be trusted to aggressively report on him? #DumpTump https://t.c
TweeetBug||0.2023|0.094|0.779|0.127|RT @GoAngelo: NBC has a financial stake in Trump's reputation. How can they be trusted to aggressively report on him? #DumpTump https://t.c
sarahblash1|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
RWNemanich|richardwolffedc|0.6369|0.0|0.785|0.215|"RT @richardwolffedc: You know, Im, like, a smart person,"" Trump tells Fox, explaining why he doesn't need intel briefings. While also pro"
