User|Original_User/Web|Compound|Negative|Neutral|Positive|Tweet
bikerbd|ColorMeRed|-0.4404|0.163|0.837|0.0|RT @ColorMeRed: Obama has no clueing  what he's accusing Russia of.. Obama has interfered with every election from Canada to Egypt... what
BillBartosik|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
adirado29|yahoo|0.0|0.0|1.0|0.0|Trump on Russia meddling in US election: 'I don't believe it' #MAGA..  https://t.co/6NYEZg1L3Y
JJFan18|MarkBrewerDems|-0.3612|0.102|0.898|0.0|RT @MarkBrewerDems: Time for reform: the legacy of @migop @MichSoS Ruth Johnson is the mess of an election system the recount revealed http
ghostwrittn|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
mommysquared|luna_sea|-0.34|0.118|0.882|0.0|"RT @luna_sea: Bipartisan group of senators say reports on Russia cyberattacks to influence election should ""alarm every American"" https://t"
mommysquared||-0.34|0.118|0.882|0.0|"RT @luna_sea: Bipartisan group of senators say reports on Russia cyberattacks to influence election should ""alarm every American"" https://t"
COBYKOEHL|NewCenturyTimes|-0.4019|0.137|0.863|0.0|RT @NewCenturyTimes: Russia Reveals Real Reason Putin Got Involved In Election; Will Piss Off Every Person https://t.co/luVrucmPbq https:/
COBYKOEHL|newcenturytimes|-0.4019|0.137|0.863|0.0|RT @NewCenturyTimes: Russia Reveals Real Reason Putin Got Involved In Election; Will Piss Off Every Person https://t.co/luVrucmPbq https:/
rememberangel00|markknoller|-0.3818|0.12|0.88|0.0|RT @markknoller: Leading network evening newscasts: CBS: Russian interference in US election?; ABC/NBC: Arctic snow and temps slam parts of
tombstone19391|schober_lisa|-0.4404|0.127|0.873|0.0|@schober_lisa @Reuters Tell me did you ask for the same thing about Hillary when she was such a train wreck through https://t.co/jzJcLfxE73
tombstone19391|twitter|-0.4404|0.127|0.873|0.0|@schober_lisa @Reuters Tell me did you ask for the same thing about Hillary when she was such a train wreck through https://t.co/jzJcLfxE73
RanttNews|casatino|-0.1027|0.097|0.903|0.0|RT @casatino: FBI: sends vague letter; actually nothingMSM: *quivers*CIA: confirms Russia interfered w/electionMSM: \_()_/https://
Eonkidz|RealAlexJones|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
Eonkidz|infowars|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
JJl500|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
Rutherfo1Melody|Green_Footballs|0.25|0.1|0.72|0.18|RT @Green_Footballs: One thing was confirmed beyond any doubt in this election: the Republican Party is just fine with white supremacism.
silentkpants|timcarvell|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
silentkpants|freep|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
asribera|UnhingedBekah|0.5046|0.0|0.86|0.14|RT @UnhingedBekah: I thought since after the results of this election anyone can be president so heres my acceptance speech @ddlovato @noma
HollieEnnissPoe|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
KenYounos|CarmineZozzora|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
KenYounos|t|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
sandlorn|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
thinkkimthink|Amy_Siskind|-0.2023|0.133|0.766|0.101|"RT @Amy_Siskind: It seems like Friday's outrage about the CIA Report and Russia's infiltrating our election, has simmered down to a whimper"
timmcdaniels|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Tabitha__Lily|RichardGrenell|0.0|0.0|1.0|0.0|"RT @RichardGrenell: Tip for @RyanLizza: If US had evidence that the Russian Government interfered with our election, we would see multiple"
denny_inspace|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
jmcrtc1|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
jmcrtc1|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
LaVerneWright13|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
LaVerneWright13|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
gamecat|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
twagz20|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
twagz20|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
PDBax|NormEisen|0.2211|0.156|0.693|0.151|@NormEisen He won election despite xenophobia. Just because people are concerned w business conflicts doesn't mean they don't want him POTUS
mchwllms5|nytimes|0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
mchwllms5||0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
valeriekeefe|iCounterSpin|0.0|0.0|1.0|0.0|"RT @iCounterSpin: If Russian's are the cause of the election, does that mean folks will lay off Berner's, Greens and Millennials now?"
dadavies|timoreilly|0.7845|0.0|0.635|0.365|"RT @timoreilly: A wonderful proposal for strengthening the civic  fabric of society, from @ericpliu. https://t.co/pFYJSgnWAC"
dadavies|theatlantic|0.7845|0.0|0.635|0.365|"RT @timoreilly: A wonderful proposal for strengthening the civic  fabric of society, from @ericpliu. https://t.co/pFYJSgnWAC"
DWGreviews|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Plantflowes|aliasvaughn|-0.2732|0.126|0.795|0.079|RT @aliasvaughn: 10. #AuditTheVote people told you straight the day after election that Russian hackers were attacking US on election night.
Shalom555222|true_pundit|-0.6124|0.318|0.547|0.135|RT @true_pundit: BuzzFeed Caught Citing Fake Data In Its Fake News Won The Election For Trump Argument  AGAIN #FakeNewshttps://t.co/mY
JPKC|socialmediatoday|0.0|0.0|1.0|0.0|How the 2016 US Presidential Election Will #socialmedia https://t.co/AS2qYrkDCz https://t.co/MVKtMnIDKE
DrSoup34|smotus|0.3164|0.144|0.642|0.214|"RT @smotus: ""Happy holidays.""""WE'RE UNDER ATTACK!""""Russia hacked our election.""""Meh, this happens all the time."""
_kaitlin_s|smotus|0.3164|0.144|0.642|0.214|"RT @smotus: ""Happy holidays.""""WE'RE UNDER ATTACK!""""Russia hacked our election.""""Meh, this happens all the time."""
Yemayah777|TazKHC|0.2924|0.0|0.902|0.098|RT @TazKHC: A bi-partisan group is challenging Trump's denial of Russian hacking in our election! Trump continuing to discredit the CIA! Lo
baloo035|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
baloo035|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
YvetteKopp|Ziggy_Daddy|0.8126|0.0|0.714|0.286|RT @Ziggy_Daddy: I never thought I'd live to see the day when Russia interferes with our election to help Trump win and Americans are okay
ParisNeully|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
complainster|aliasvaughn|-0.3348|0.117|0.883|0.0|RT @aliasvaughn: @davebernstein DOJ numbers here . CALL!!! Demand full investigation on Russia hacks/comey/trump AND audit and redo of elec
mikemovie|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
Ruth_elsesser|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
fruitfriend|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
anamerican397|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
cecilia_c_chung|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
heatherdean71|Neighbors4Hill|0.0|0.0|1.0|0.0|RT @Neighbors4Hill: Call Mitch McConnell 202-224-2541 to ask him why he kept us in the dark about foreign interference in our election
tony_thetruth|1Marchella|-0.1531|0.078|0.922|0.0|"RT @1Marchella: ""We've got no evidence that #RussianHackers influenced the election, but we're going to report they did anyway"" https://t.c"
tony_thetruth||-0.1531|0.078|0.922|0.0|"RT @1Marchella: ""We've got no evidence that #RussianHackers influenced the election, but we're going to report they did anyway"" https://t.c"
grumpee_mike|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
Dimipace|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Dimipace||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
CPTsopiens|seanmdav|-0.8176|0.292|0.664|0.043|"RT @seanmdav: Is the NFL still blaming the election for this, or have they moved on to another stupid excuse no one buys? https://t.co/OXga"
CPTsopiens|t|-0.8176|0.292|0.664|0.043|"RT @seanmdav: Is the NFL still blaming the election for this, or have they moved on to another stupid excuse no one buys? https://t.co/OXga"
CAGoldenBear|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
DiggleLynn|TrumpsNewsDaily|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
DiggleLynn|yahoo|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
sabretoothsdrum|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Beverly86418528|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
DarienBresee|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
DarienBresee|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
DragoEldur|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
AndrewKayNZ|twitter|0.3412|0.0|0.893|0.107|"You won't have to worry about the next election, the way labour is polling, you'll probably be rolled by then. https://t.co/RYgToCi1yt"
Ish|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
RMB_Investor|rmbinvestor|0.0|0.0|1.0|0.0|"Ld 's Hk Chief Executive Says Not To Seek Re Election  : https://t.co/4zGz9NLRb6 ,"
HonestPolitics7|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Awtcaribbean|politico|0.0|0.0|1.0|0.0|Obama orders 'deep dive' of election-related hacking https://t.co/DudYfoiTB3
AndreFrato|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Karen6349|DavidAFrench|-0.3612|0.122|0.878|0.0|RT @DavidAFrench: What's the argument against a bipartisan investigation of Russian efforts to disrupt and/or influence the election? Is th
MtRushmore2016|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Benst90|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
BudtPert|greenhousenyt|-0.0516|0.11|0.787|0.102|"RT @greenhousenyt: ""The fact that 59% of the vote-counting machines in Detroit all broke on Nov. 8 stands out as a stunning developmnt"" htt"
AbhijitVaidya|heytal|-0.3182|0.18|0.735|0.086|"@heytal no. Visited Chinchwad yesterday. There were a lot of those. In pune, no of hoardings are increased in general, considering election"
BonnieSue05060|summerbrennan|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
BonnieSue05060|t|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
PAposter|palmerreport|-0.4215|0.157|0.843|0.0|Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/4mhK9gYmIS
Angelmdunn1961|PrisonPlanet|-0.5106|0.191|0.809|0.0|"RT @PrisonPlanet: Post election riots: FAILED.Jill Stein recount: FAILED.Intimidation of EC members: FAILED.""Fake news"": FAILED.""Russia"
angelfrmcanada|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
angelfrmcanada|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
parandersj|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
parandersj||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
Winston_Truth|Neighbors4Hill|0.0|0.0|1.0|0.0|RT @Neighbors4Hill: Call Mitch McConnell 202-224-2541 to ask him why he kept us in the dark about foreign interference in our election
Tabitha__Lily|SaysSimonson|-0.4588|0.13|0.87|0.0|RT @SaysSimonson: @RichardGrenell @RyanLizza the people attacking trump for the intel briefings are the same people who reported on an elec
tardiskitten|greenhousenyt|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
tardiskitten|t|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
jackthecat111|timcarvell|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
jackthecat111|freep|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
pandagabe|CEDADebate|0.7345|0.0|0.754|0.246|"RT @CEDADebate: The election results are in, thank you to everyone who ran and congrats to everyone who was elected!... https://t.co/nh5AFX"
pandagabe|t|0.7345|0.0|0.754|0.246|"RT @CEDADebate: The election results are in, thank you to everyone who ran and congrats to everyone who was elected!... https://t.co/nh5AFX"
TINTofPBC|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
CynicalParadox|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
KattNasty|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
sanjerina|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
maryjane0250|Moo57556470|-0.5994|0.151|0.849|0.0|"RT @Moo57556470:  Isn't the #RussianHacking to compromise our election an act of cyber war? Is PEOTUS, Congress &amp; Comey's FBI on our si"
linda_wed1|PolticsNewz|-0.4404|0.146|0.854|0.0|RT @PolticsNewz: Sen. Mitch McConnell needs to answer for his role covering up Russian election attacks https://t.co/p083ik11O3 https://t.c
linda_wed1|route|-0.4404|0.146|0.854|0.0|RT @PolticsNewz: Sen. Mitch McConnell needs to answer for his role covering up Russian election attacks https://t.co/p083ik11O3 https://t.c
D_TownFan|ed_hooley|-0.5754|0.157|0.843|0.0|RT @ed_hooley: JOHN MCCAIN: RUSSIA HACKED OUR ELECTION! MCCAIN IS BOUGHT &amp; SOLD BY GEORGE SORO'S #McCain #JohnMcCain #Arizona #teaparty htt
Mannyratback1|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Our favourite #FakeNews of the 2016 election https://t.co/Onm82JGBbn
Mannyratback1|twitter|0.0|0.0|1.0|0.0|RT @wikileaks: Our favourite #FakeNews of the 2016 election https://t.co/Onm82JGBbn
Iangroome|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
CaridadDorado|nytimes|0.4767|0.0|0.853|0.147|RT @nytimes: Breaking News: President Obama orders intelligence agencies to report on Russian efforts to influence 2016 election https://t.
CaridadDorado||0.4767|0.0|0.853|0.147|RT @nytimes: Breaking News: President Obama orders intelligence agencies to report on Russian efforts to influence 2016 election https://t.
SabraJewell|mhmck|-0.3818|0.12|0.88|0.0|"@mhmck @M5B1tch Obama declare State of emergency, stays in office till 2018 midterms, New GOP candidate, redo the National Election"
Hasfot7|ABC|0.0|0.0|1.0|0.0|RT @ABC: NEW: Bipartisan group of senators release joint statement calling for examination of reports of Russian interference in 2016 US el
HH75876116|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
BigTimeCarly|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
piyamoda|sygebowyf|0.0|0.0|1.0|0.0|RT @sygebowyf: WASHINGTON  An extraordinary breach has emerged between President-elect Donald  https://t.co/0Fhtmj0P7f
piyamoda|nytimes|0.0|0.0|1.0|0.0|RT @sygebowyf: WASHINGTON  An extraordinary breach has emerged between President-elect Donald  https://t.co/0Fhtmj0P7f
jbtcarolina|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
MyNameIsSergius|mtracey|-0.2263|0.102|0.837|0.06|@mtracey With no proof of hacking during the election they want a new vote eh? Here's my answer to them - https://t.co/sIAr4UCmqD
MyNameIsSergius|twitter|-0.2263|0.102|0.837|0.06|@mtracey With no proof of hacking during the election they want a new vote eh? Here's my answer to them - https://t.co/sIAr4UCmqD
SissyWarf|WFMY|0.0|0.0|1.0|0.0|RT @WFMY: Trump dismisses allegations of Russian election tampering https://t.co/BrqMbgYJq7 https://t.co/goZW8NiGD0
SissyWarf|wfmynews2|0.0|0.0|1.0|0.0|RT @WFMY: Trump dismisses allegations of Russian election tampering https://t.co/BrqMbgYJq7 https://t.co/goZW8NiGD0
ShitCanUrCoach|realDonaldTrump|-0.7003|0.254|0.746|0.0|"@realDonaldTrump the dems would have chose some Berkeley dumbass theoretitian, with no experience... that worked for obama, election showed"
DonnyDidntDoIt|medium|-0.3736|0.146|0.854|0.0|"Was this the objective? #republicans stop #merrickgarland, #donaldtrump deal w/ #russia &amp; #putin hacks election? https://t.co/JZntohKemP"
terebifunhouse|timcarvell|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
terebifunhouse|freep|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
vela_mary|JuddLegum|0.4404|0.0|0.847|0.153|RT @JuddLegum: Updated list of GOP members supporting investigation into Russian interference w/prez electionSen GrahamSen McCainSen Co
Discoexpress|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: New SMS records show Assange was framed by police in 1st sex case: https://t.co/MqwZAvH0va and in 2nd case: https://t.co/OPC
Discoexpress|justice4assange|0.0|0.0|1.0|0.0|RT @wikileaks: New SMS records show Assange was framed by police in 1st sex case: https://t.co/MqwZAvH0va and in 2nd case: https://t.co/OPC
BelkysSpainUSA|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
suicide_romance|casatino|-0.1027|0.097|0.903|0.0|RT @casatino: FBI: sends vague letter; actually nothingMSM: *quivers*CIA: confirms Russia interfered w/electionMSM: \_()_/https://
mymeraki1|ArvindKejriwal|-0.296|0.087|0.913|0.0|@ArvindKejriwal all time u putting aligation on pm that he stop me working in Delhi and I think u'll be say same lines after Punjab election
scudderplus|johnmccain2016|-0.5106|0.142|0.858|0.0|@johnmccain2016 your outrage over the Russian hack would have carried more weight had you shown a spine against Trump during the election.
ActorAaronBooth|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
ActorAaronBooth|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
ItsaVapeThang|HEROESvape|0.296|0.0|0.864|0.136|RT @HEROESvape: Im busy creating enough white clouds to signal the election of a new pope.
marcirish|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
Badgersbane|birbigs|-0.0387|0.05|0.95|0.0|RT @birbigs: There's evidence that Russia swayed the U.S. election &amp; we're supposed to NOT talk about it constantly? I'm sorry but that's u
laun|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
aaron_rva|YouTube|0.0|0.0|1.0|0.0|I added a video to a @YouTube playlist https://t.co/RcFJO6qsx0 MSNBC Election Night 2016 Full Coverage 2/3 (No Commercials)
aaron_rva|youtube|0.0|0.0|1.0|0.0|I added a video to a @YouTube playlist https://t.co/RcFJO6qsx0 MSNBC Election Night 2016 Full Coverage 2/3 (No Commercials)
IamSilverPeace|MadJewessWoman|0.0|0.0|1.0|0.0|"RT @MadJewessWoman: .@realDonaldTrumpINVESTIGATE @SenJohnMcCain 4 overthrowing #Ukraine govt, influencing election in #KIEV, 2013-14http"
DawnQuesarrah|bonita_jay1|0.0772|0.0|0.936|0.064|RT @bonita_jay1: @kirangkaur @aliasvaughn There is a petition to indicate that this is precisely what US citizens want to happen: https://t
DawnQuesarrah||0.0772|0.0|0.936|0.064|RT @bonita_jay1: @kirangkaur @aliasvaughn There is a petition to indicate that this is precisely what US citizens want to happen: https://t
StrellcZeneli|youtube|-0.2023|0.153|0.847|0.0|Islamic scholar Imran Hosein: Trump's election may have postponed nuclea... https://t.co/gktcxfhHVe
SamanthaMakoski|twitter|-0.3182|0.247|0.753|0.0|This election is making for odd bedfellows. https://t.co/3vX9QPVmru
annetteKwest|TuckerCarlson|0.5859|0.0|0.798|0.202|"RT @TuckerCarlson: President-elect @realDonaldTrump to protester: The election ended 3 weeks ago, darling TCT #Tucker @FoxNews https://t"
annetteKwest||0.5859|0.0|0.798|0.202|"RT @TuckerCarlson: President-elect @realDonaldTrump to protester: The election ended 3 weeks ago, darling TCT #Tucker @FoxNews https://t"
IBDeb2|latimes|0.0|0.0|1.0|0.0|This shouldn't be a partisan issue. It is an American issue. Disturbing/telling thatTrump doesn't see it that way    https://t.co/Uz5lciHGBU
jmarong69|Engelkes|0.7003|0.084|0.649|0.267|RT @Engelkes: No sitting Supreme Court in #Gambia. Current chief justice is Nigerian. 4 other judges to be hired https://t.co/DonEFu2Orz vi
jmarong69|reuters|0.7003|0.084|0.649|0.267|RT @Engelkes: No sitting Supreme Court in #Gambia. Current chief justice is Nigerian. 4 other judges to be hired https://t.co/DonEFu2Orz vi
VickyDurieux|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
VickyDurieux||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
LiMystery|realDonaldTrump|0.5719|0.0|0.837|0.163|"If #RussiaHacking results in a new election and @realDonaldTrump wins AGAIN, facts haven't changed,so why not call for ANOTHER new election?"
jackthecat111|timcarvell|-0.34|0.107|0.893|0.0|RT @timcarvell: @markoff The election official goes on to say that not all precincts would necessarily be excluded for this reason.
lorax58|MrJamesonNeat|-0.6597|0.231|0.769|0.0|RT @MrJamesonNeat: In states where election fraud seems rampant lawsuits should be filed to disqualify Trump electors @tribelaw @lessig htt
michaels_leigh|iveygirl08|0.0|0.0|1.0|0.0|RT @iveygirl08: Latest Election Results: Congressman Calls On Elec... https://t.co/ogI6BIHWxp
michaels_leigh|topbuzzapp|0.0|0.0|1.0|0.0|RT @iveygirl08: Latest Election Results: Congressman Calls On Elec... https://t.co/ogI6BIHWxp
BossClaw|SafeWordApples|-0.8271|0.303|0.697|0.0|RT @SafeWordApples: Russia hacked the election is 2016's the dog ate my homework. One of the stupidest excuses for losing an election. #Rus
JudyThompson13|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
NYtitanic1999|UKChange|0.0|0.0|1.0|0.0|President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/ifEZvwtJgx via @UKChange
NYtitanic1999|linkis|0.0|0.0|1.0|0.0|President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/ifEZvwtJgx via @UKChange
fairservice_3|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
ValRayOSunshine|Vote_American|-0.6407|0.225|0.775|0.0|RT @Vote_American: Didn't United States (Obama) meddled in Israeli Last Election by funding efforts to Unseat Netanyahu? Obama hates him. O
misssqueakums|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
suemagic|M|0.0|0.0|1.0|0.0|Rep. John Lewis has submitted a bill to Congress authorizing a 2nd National Election. call reps (202) 224-3121 https://t.co/sxJeXjBkfA
DSTrey5|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
TeamTrumpTeX|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
MacneilAl|michaelianblack|0.4404|0.0|0.828|0.172|@michaelianblack Just look at your investment performance since election; that'll make you feel better #trumpeconomy
chris_wtu|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
MikeJr8282|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
M_CollinsDesign|HouseofCards|-0.0429|0.104|0.798|0.098|America was so impatient for new seasons of @HouseofCards &amp; @VeepHBO that we made the 2016 election to keep us entertained in the meantime.
fscheune1|nytimes|0.0|0.0|1.0|0.0|https://t.co/HFKrlC91MQ
sarahrivell|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
sarahrivell|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
mountainman7|_Makada_|-0.296|0.115|0.826|0.06|"RT @_Makada_: President-Elect Trump: It's ridiculous to say Russia intervened in the election, I think it's just another excuse. We had a m"
morgan_blade|maddow|-0.1531|0.18|0.699|0.121|"RT @maddow: We now have high confidence they hacked the DNC and RNC, and conspicuously released no documents from the RNC https://t.co/Ue"
morgan_blade|t|-0.1531|0.18|0.699|0.121|"RT @maddow: We now have high confidence they hacked the DNC and RNC, and conspicuously released no documents from the RNC https://t.co/Ue"
mgyousey|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
jevans15|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
heinemannp|sacca|0.6369|0.088|0.654|0.258|RT @sacca: On @NPR I shared why tech leaders who go to Trump Tower will get played and also lose the respect of employees. https://t.co/XGA
heinemannp|t|0.6369|0.088|0.654|0.258|RT @sacca: On @NPR I shared why tech leaders who go to Trump Tower will get played and also lose the respect of employees. https://t.co/XGA
abs_tellthetale|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
jenscorpio83|Neighbors4Hill|0.0|0.0|1.0|0.0|RT @Neighbors4Hill: Call Mitch McConnell 202-224-2541 to ask him why he kept us in the dark about foreign interference in our election
mariecasey1|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
tsubi|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
newacademic|mtracey|-0.25|0.095|0.905|0.0|"RT @mtracey: Dems' post-election lunacy closely resembles GOP birtherism, except in this case the paranoia is far more mainstream https://t"
newacademic||-0.25|0.095|0.905|0.0|"RT @mtracey: Dems' post-election lunacy closely resembles GOP birtherism, except in this case the paranoia is far more mainstream https://t"
rogiloc|Karin_Winski|-0.4574|0.272|0.728|0.0|RT @Karin_Winski: Damn right! #NotMyComrade #TreasonousGOP #riggedelection #RevoteNow https://t.co/cEYLc8O6G5
rogiloc|politicususa|-0.4574|0.272|0.728|0.0|RT @Karin_Winski: Damn right! #NotMyComrade #TreasonousGOP #riggedelection #RevoteNow https://t.co/cEYLc8O6G5
Sharonnemesio|heatstreet|0.4588|0.0|0.864|0.136|"@heatstreet The rise of unelected, actors, 'celebrities', journalists trying to dictate to the people.   Grateful for the election of Trump"
TeckieGirl|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
SharonS72105601|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
WildlifeNRacing|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
TurnTNBlue|bannerite|-0.1027|0.1|0.815|0.085|"RT @bannerite: Mark my word, @CIA knows for sure that Russia hacked our election. But they can't reveal sources without putting them at ris"
SpazP|randysusanmeyer|0.0|0.0|1.0|0.0|RT @randysusanmeyer: Weigh in on Fox News poll!! Q: Should the U.S. investigate allegations of Russian interference in the election?https:/
SpazP||0.0|0.0|1.0|0.0|RT @randysusanmeyer: Weigh in on Fox News poll!! Q: Should the U.S. investigate allegations of Russian interference in the election?https:/
crawforddel3|randyprine|0.0|0.0|1.0|0.0|RT @randyprine: So Comey does THIS knowing the CIA has evidence that Russia was ALREADY tampering with the balance of the election. What a
aliasvaughn|summerbrennan|-0.4767|0.163|0.837|0.0|"RT @summerbrennan: As I've said before, I called McCain and Graham offices multiple times in tears right after the election and they are no"
markvukovic|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
markvukovic|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
danielj_horn|DaniSButcher|0.6369|0.0|0.769|0.231|RT @DaniSButcher: The best part about liberals saying Russia interfered with our election is: https://t.co/5rtYqDob7D
danielj_horn|twitter|0.6369|0.0|0.769|0.231|RT @DaniSButcher: The best part about liberals saying Russia interfered with our election is: https://t.co/5rtYqDob7D
Marypat714|neilpX|-0.5423|0.17|0.83|0.0|"RT @neilpX: If McCain and Graham are able to expose the treason promulgated in the election, they will deserve to be heralded as American h"
wellfedred|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
wellfedred|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
AJVicens|rickhasen|-0.0772|0.08|0.92|0.0|RT @rickhasen: #ELB; Sorry But Alleged Russian Influence in Presidential Election Wont Lead to a Do-Over https://t.co/qRyNjiCXmh
AJVicens|electionlawblog|-0.0772|0.08|0.92|0.0|RT @rickhasen: #ELB; Sorry But Alleged Russian Influence in Presidential Election Wont Lead to a Do-Over https://t.co/qRyNjiCXmh
annfinster|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
annfinster|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Coquietchat|washingtonpost|0.7579|0.0|0.683|0.317|The CIA has concluded that Russia intervened to help Trump win the US election. https://t.co/ieRdgCOq1M https://t.co/ZyVGQtMTVe
qkode|qkode|0.5423|0.0|0.774|0.226|"RT @qkode: Optimism on economy, stocks surges since Trump election: CNBC survey.. https://t.co/INMW9raLI9"
qkode|cnbc|0.5423|0.0|0.774|0.226|"RT @qkode: Optimism on economy, stocks surges since Trump election: CNBC survey.. https://t.co/INMW9raLI9"
RealAndyPanda|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
StefanHayden|PattyMurray|0.3182|0.0|0.905|0.095|RT @PattyMurray: An investigation must begin as soon as possible on any evidence Russia actively worked to hijack our election &amp; elect Dona
ReallyDontTrump|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
Donna_DHKBB|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
AliciaHallCO|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
JulieForeman16|duanecaldwell|0.4019|0.0|0.881|0.119|RT @duanecaldwell: Why is Obama now interested in Russian interference in the election?He sat around months before it and did nothing.htt
GadflyQuebec|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
maturewisdom|ECpetition|0.0|0.0|1.0|0.0|RT @ECpetition: https://t.co/6SdQhpNUQv
maturewisdom|nytimes|0.0|0.0|1.0|0.0|RT @ECpetition: https://t.co/6SdQhpNUQv
bhmoll5000|twitter|-0.2247|0.189|0.7|0.111|"I think I can help w the whole ""who really hacked the election &amp; allowed Putins surgically augmented cock to be thr https://t.co/ZUqrzbXy55"
suicide_romance|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
wolverinelmj|danversohara|0.0|0.0|1.0|0.0|RT @danversohara: Everyone around me: the election is over get over itMe: https://t.co/ykfoZyr5k2
wolverinelmj|twitter|0.0|0.0|1.0|0.0|RT @danversohara: Everyone around me: the election is over get over itMe: https://t.co/ykfoZyr5k2
JkFlower60|JasonKander|-0.6597|0.213|0.787|0.0|"RT @JasonKander: If we ignore Russian espionage in our election, we embolden other foreign powers to launch similar attacks on every aspect"
LaCina52|cdelbrocco|-0.6342|0.188|0.812|0.0|RT @cdelbrocco: He's a fucking liar!! Trump: It's 'Ridiculous' To Think Russia Intervened In The Election On My Behalf  https://t.co/hI0W
LaCina52|t|-0.6342|0.188|0.812|0.0|RT @cdelbrocco: He's a fucking liar!! Trump: It's 'Ridiculous' To Think Russia Intervened In The Election On My Behalf  https://t.co/hI0W
kvg1988|JanJohnsonFL|-0.5707|0.257|0.644|0.099|@JanJohnsonFL @kurteichenwald libtards were sure about the election... the recounts... and now the Russian hacker conspiracy! They're lost.
NedSparks|BrendanNyhan|-0.4659|0.169|0.787|0.043|"RT @BrendanNyhan: Seeing people dismiss as silly conspiracy talk, but far more serious. Potential Dep SOS suggesting Obama used IC in a dom"
JeffersonsNotes|westernlvr|0.0|0.0|1.0|0.0|@westernlvr @WalshFreedom @NBCNews These people are just reporting what the Russians said!!!! Here's Fortune.https://t.co/QHYQdHA3Ac
ElenaSryva|kurteichenwald|-0.2382|0.22|0.67|0.11|"RT @kurteichenwald: No offense, @chucktodd, but when u say no one was sure Russia behind hack pre-election, shows u need to read more. http"
mbrobison|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
mbrobison||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
luna_sea|npr|-0.34|0.13|0.87|0.0|"Bipartisan group of senators say reports on Russia cyberattacks to influence election should ""alarm every American"" https://t.co/2ce7PoYTR5"
donalds_dad|twitter|-0.1027|0.076|0.924|0.0|#TeamTrump challenged the veracity of US intel that Russia influenced #election for #Trump. Not what #Russia intel https://t.co/wi7NKMOt6m
katomart|MarkDice|0.0|0.183|0.633|0.183|RT @MarkDice: Stop.  You idiots failed in all your predictions about the election. Just accept that Trump is better in every way. https://t
katomart||0.0|0.183|0.633|0.183|RT @MarkDice: Stop.  You idiots failed in all your predictions about the election. Just accept that Trump is better in every way. https://t
karenkho|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
MikeJC12019|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
crankonosborn|abermans|-0.3802|0.126|0.874|0.0|RT @abermans: 2/2017 #Election?Come what #may wants:More #Brexit delay and more tory power.Only she will get mass #UKIP upvote!https://
crankonosborn||-0.3802|0.126|0.874|0.0|RT @abermans: 2/2017 #Election?Come what #may wants:More #Brexit delay and more tory power.Only she will get mass #UKIP upvote!https://
RB98SS|steph93065|-0.296|0.104|0.896|0.0|@steph93065 They knew it'd take 12yrs to fundamental Transform Amer an without HRC their screwed.They'll do anything to undermine election.
VLaw09|jameshamblin|0.0|0.0|1.0|0.0|RT @jameshamblin: So people believe a pizza place is a government sex ring but fancy themselves too savvy to look into Russian election int
vancetran|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
scandalholic|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
scandalholic||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
NickEKnockers|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
sethsoren|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
AltRockAddict|Holbornlolz|-0.6705|0.231|0.684|0.085|RT @Holbornlolz: People who killed 100's of 1000's to ensure regime change all over the M. East are upset that Russia may have interfered i
LegalForTrump|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
siempreuntigre|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
CerridwenF|facebook|0.0|0.0|1.0|0.0|Keep throwing it all against the wall--maybe something will stick...Russian interference in our election makes... https://t.co/PLyZZzWdWP
SheriHerman10|Counter_info|-0.4019|0.231|0.769|0.0|@Counter_info Its utter BS that Russia hacked the US election.
ciaobella50|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
runnin5|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
tom_klem|GeorgeTakei|0.34|0.0|0.902|0.098|"RT @GeorgeTakei: If there was interference on the play, you don't count the touchdown. Russia meddled in our election, says the CIA. Electo"
gibson_marianne|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: Also, there must be investigation of Comey @FBI. That he could know this &amp; decide to break all history to interfere w/"
cakehler|RepublicanChick|-0.1779|0.082|0.918|0.0|"RT @RepublicanChick: Liberals are accusing Russia of influencing the election. At the same time, liberals enabled citizens of other countri"
d10r10_jeremy|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: What if the election hadn't been hacked?What if Hillary hadn't stole the nomination?What if Obama hadn't given rise to
Daniel_Ross622|DavidAFrench|-0.3612|0.122|0.878|0.0|RT @DavidAFrench: What's the argument against a bipartisan investigation of Russian efforts to disrupt and/or influence the election? Is th
Jordan_Milam|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
slidewinding|jahimes|0.6375|0.0|0.754|0.246|RT @jahimes: @GoodJobGuru @PoliticalLine Yes. The election is over. But the electoral college has not met. So no President has been legally
verna_williams|birbigs|-0.0387|0.05|0.95|0.0|RT @birbigs: There's evidence that Russia swayed the U.S. election &amp; we're supposed to NOT talk about it constantly? I'm sorry but that's u
CintiNative|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
CintiNative|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Robertvest1Vest|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
Grumpy_Ol_Me|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ftvoc|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
heathergilding|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
alitaleader|twitter|-0.3612|0.156|0.844|0.0|"These boots are made for walking, we need to walk right to DC and protest the election and demand a revote.Thanks, https://t.co/NrVE96SqND"
Searching4Par|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
vmsre|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
LizKennedy_|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
LizKennedy_||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
benfinzel|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
eclubproject|mashable|0.0|0.0|1.0|0.0|RT @mashable: The one social platform actually taking action ahead of Trump's America https://t.co/4Q3d2SnM5G https://t.co/41TlUUVzx2
eclubproject|mashable|0.0|0.0|1.0|0.0|RT @mashable: The one social platform actually taking action ahead of Trump's America https://t.co/4Q3d2SnM5G https://t.co/41TlUUVzx2
Kane_Says405|Shoq|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
Kane_Says405|t|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
Wadatahmydamie|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Mannyratback1|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Mannyratback1|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
tpinklittle|DecksDarkAlien|0.0|0.0|1.0|0.0|"RT @DecksDarkAlien: So, the story begins in WaPo as a ""he said she said"" report &amp; now, media everywhere reports it as a CIA report? https:/"
tpinklittle||0.0|0.0|1.0|0.0|"RT @DecksDarkAlien: So, the story begins in WaPo as a ""he said she said"" report &amp; now, media everywhere reports it as a CIA report? https:/"
BevPerryMusic|amjoyshow|0.0|0.0|1.0|0.0|"RT @amjoyshow: Will Donald Trump's election empower African ""strongmen"" dictatorial rulers? Our panel goes in #AMJoy https://t.co/AddWC2TuYB"
BevPerryMusic|twitter|0.0|0.0|1.0|0.0|"RT @amjoyshow: Will Donald Trump's election empower African ""strongmen"" dictatorial rulers? Our panel goes in #AMJoy https://t.co/AddWC2TuYB"
Zoraida12098036|DailyNewsBin|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
Zoraida12098036|palmerreport|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
LuckyDuckyToo|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
Lazer_Mondass|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
Lazer_Mondass|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
Ldyforce6|AlexUSA1956|-0.0516|0.162|0.684|0.154|"RT @AlexUSA1956: Supreme Court: Election Can Be Invalidated Due To Massive Fraud, Install Opponent (DETAILS) https://t.co/WEH9OdQIX6 via @B"
Ldyforce6|bipartisanreport|-0.0516|0.162|0.684|0.154|"RT @AlexUSA1956: Supreme Court: Election Can Be Invalidated Due To Massive Fraud, Install Opponent (DETAILS) https://t.co/WEH9OdQIX6 via @B"
realNiggaTrump|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
PDI_Proyectos|washingtonpost|0.7579|0.0|0.667|0.333|The CIA has concluded that Russia intervened to help Trump win the US election. https://t.co/yRwoo2Qq2p
slickvolt|washingtonpost|0.1027|0.117|0.745|0.138|@washingtonpost @ABC @CBSNews @CNN @FoxNews @NBCNews @MSNBC UNAMERICAN Democrat politicians refuse to accept results of election...LIARS
luvthmgators|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
lkaiser8|colinjones|0.3182|0.116|0.677|0.207|"RT @colinjones: You know, Im, like, a smart person. - Trump on criticism of his refusal of more regular intel briefings https://t.co/aGd"
lkaiser8|t|0.3182|0.116|0.677|0.207|"RT @colinjones: You know, Im, like, a smart person. - Trump on criticism of his refusal of more regular intel briefings https://t.co/aGd"
ElizbethLManess|WeNeedTrump|-0.4522|0.129|0.871|0.0|"RT @WeNeedTrump: So the left cries about Russia allegedly interfering with our election. Yet, millions were donated to the Clinton Foundati"
issuemaverick|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
MissLin68640163|JYSexton|-0.7003|0.264|0.652|0.084|RT @JYSexton: And for what? The election of a man who disgusts them and makes a mockery of their party. What a sad sack of shills these peo
beatthebrain|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
LEngelhorn|aliasvaughn|-0.3597|0.102|0.898|0.0|"RT @aliasvaughn: 9. So stop trying with ""oh they just ""tried to influence"" the election"" and start realizing that what we're dealing with i"
TheDon2174|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
NicoDeWitty|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
TimLimDC|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
CCFPHD|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
CCFPHD||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
RLSRUSSIANNEWS|theguardian|0.0|0.0|1.0|0.0|Donald Trump says CIA charge Russia influenced election is 'ridiculous' - The Guardian https://t.co/1vXW7UbF3J
RichardCalahan|JohnWDean|0.0|0.0|1.0|0.0|RT @JohnWDean: The intel report on Russia's role in the 2016 election must be available for all electors before the electoral college meets
HankPettit|RepublicanChick|-0.1779|0.082|0.918|0.0|"RT @RepublicanChick: Liberals are accusing Russia of influencing the election. At the same time, liberals enabled citizens of other countri"
wigbayer|LeahR77|0.1531|0.11|0.758|0.133|RT @LeahR77: Lets Talk Foreign Govts Influencing An Election &amp; Bonus Getting Uranium &amp; Weapons Deals From SOS HRC For #FakeNews #Russians
Cwmateo|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
hopefor_america|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
iantothemax|2dJazz|0.7845|0.0|0.685|0.315|RT @2dJazz: Arc System Works Awards 2016 election results:GG: @koichinko &amp; @gou4th_fab BB: @soujif91 &amp; @MINAMI_IZANAMI Congratulations 
MelissaHoughto6|Trump4Pres0225|-0.5106|0.148|0.852|0.0|RT @Trump4Pres0225: .@POTUSwas given Morning briefs on CIA concerns with Russia involvement PRE ELECTION.  Where was the outrage THEN? http
bikerbd|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
bikerbd|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
annemelvinbloom|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
annemelvinbloom|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
edgeoforever|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: MOVING ON. The conspiratorial fever at about 108, we begin the 2016 election - AGAINST EVERYTHING HOLY - in 2015."
Dr_2A|ctalmon|0.5106|0.0|0.829|0.171|Feel free to have an alternate opinion of what hack the election means.Where is this evidence?@ctalmon @walshfreedom
OurPowderDry|davidfrum|0.0|0.0|1.0|0.0|@davidfrum Obama needs to link Russia/Trump collusion now. Friday WH news big game changer but 2 little 2 late. https://t.co/S2m37OCzm7
OurPowderDry|change|0.0|0.0|1.0|0.0|@davidfrum Obama needs to link Russia/Trump collusion now. Friday WH news big game changer but 2 little 2 late. https://t.co/S2m37OCzm7
Michael26222747|JLynn8412|-0.4588|0.188|0.735|0.077|RT @JLynn8412: @JuddLegum well @SenateMajLdr is the leader of treason as he refused to let info. out to public before election. Why would h
ParthPatel9|AoDespair|-0.3885|0.192|0.638|0.17|RT @AoDespair: Fucking hell. National health care? Response to global warming? Sending a man to Mars? We can't even run a functional electi
WinterDaisy|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
SN_Tobin|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
SN_Tobin||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Jaxon_Dillinger|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ChanCans529|EvelKnievel5|-0.2732|0.227|0.623|0.15|RT @EvelKnievel5: @Magdaletou @funder are you still sad about the election cupcake?  That was a great night watching libs cry https://t.co/
ChanCans529|t|-0.2732|0.227|0.623|0.15|RT @EvelKnievel5: @Magdaletou @funder are you still sad about the election cupcake?  That was a great night watching libs cry https://t.co/
Rudedog6557|MaydnUSA|-0.4019|0.119|0.881|0.0|"RT @MaydnUSA: When Sony was hacked, the FBI immediately produced evidence. Anyone seen any actual evidence of election hack by Russia?Did"
Robotbeat|ericgarland|0.0|0.0|1.0|0.0|"RT @ericgarland: MOVING ON. The conspiratorial fever at about 108, we begin the 2016 election - AGAINST EVERYTHING HOLY - in 2015."
atriverside|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
bulletin_world|theworldbulletin|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votescounted https://t.co/GCRwAjZ32C https://t.co/7MXSPOOhZ1
sabine_durden|wraithvenge|-0.4215|0.268|0.606|0.126|RT @wraithvenge: .@riyasharma266 Just like she abandoned them on election night when she lost https://t.co/uPKUP3NUp9
sabine_durden|twitter|-0.4215|0.268|0.606|0.126|RT @wraithvenge: .@riyasharma266 Just like she abandoned them on election night when she lost https://t.co/uPKUP3NUp9
algonzalezlu393|Pinkcloud15|0.2225|0.0|0.914|0.086|RT @Pinkcloud15: It's time 2 take our country back! Call the W H 202-456-1414 'n tell thm U want a new election done w/paper ballots! https
WandaMiller5102|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
WandaMiller5102|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
GaTo_TrenDy|twitter|0.2023|0.0|0.878|0.122|Trump faces first significant post-election pushback from Republicans over CIA report on Russia https://t.co/pgDIUVRhf4
SunnyJL52|Irwin_Elaine|0.0|0.0|1.0|0.0|RT @Irwin_Elaine: @_0HOUR1 Here's a list of all the Foreign Governments who interfered in the last Pres election. I mean... donated to the
mccay_rl|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
Real_TrumpFacts|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
hecksmaniac|2dJazz|0.7845|0.0|0.685|0.315|RT @2dJazz: Arc System Works Awards 2016 election results:GG: @koichinko &amp; @gou4th_fab BB: @soujif91 &amp; @MINAMI_IZANAMI Congratulations 
keating_eleanor|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
DeBellSar|leahmcelrath|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
DeBellSar|t|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
DrKousigan|HuffPostPol|-0.5719|0.236|0.764|0.0|RT @HuffPostPol: Bipartisan anger grows over Russian interference into U.S. election https://t.co/YOujihnfxw https://t.co/IGTG7ysCMG
DrKousigan|m|-0.5719|0.236|0.764|0.0|RT @HuffPostPol: Bipartisan anger grows over Russian interference into U.S. election https://t.co/YOujihnfxw https://t.co/IGTG7ysCMG
islamophobie2|barenakedislam|0.0|0.0|1.0|0.0|FLYING PIGS MOMENT from a far left writer at the New York Times: Election https://t.co/ik8lOh0Idu #islamofobia
dougsheridan|mtracey|0.0|0.0|1.0|0.0|"@mtracey Right, cuz ex-CIA operatives are always the last word when it comes to Presidential-election redos. #fakecnnnews"
PatLynnFor|twitchy|0.0|0.0|1.0|0.0|"McCain is a WEASEL:  Graham, McCain,Schumer and Reed release joint statement on Russian interference w/2016 election https://t.co/fynuHArbEf"
NotAmandaW|sethmoulton|0.6808|0.0|0.811|0.189|"RT @sethmoulton: Proud to see so many #MA6 constituents ready to work for change. There is so much to do, and this election was a call to a"
FWjmcg|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
FWjmcg|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Teacher4Sanders|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
RedRose3b|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
RedRose3b||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
creekbear|NarratedPOTUS|0.4019|0.139|0.623|0.238|RT @NarratedPOTUS: The President-elect of the United States asserts that there was rampant voter fraud in the election he won.
ProfTowanda|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
ProfTowanda||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
RenegadeB3|PrisonPlanet|-0.3453|0.139|0.861|0.0|RT @PrisonPlanet: Russia interfered in the election! (no evidence).LEFT FREAKS OUT.Saudi Arabia provably bankrolled Clinton's campaign.
globalissuesweb|twib|-0.4767|0.437|0.563|0.0|Nigeria: Election Suspended https://t.co/l0XBIui5XC https://t.co/Ir299AuhQa
jhanmuoz1|twitter|0.2023|0.0|0.878|0.122|Trump faces first significant post-election pushback from Republicans over CIA report on Russia https://t.co/jnwwd4HFop
Lou74inKC|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
tweeharley823|DavidYankovich|-0.296|0.109|0.891|0.0|RT @DavidYankovich: There is no Democrat/Republican side to the Russian influence in this election.You are either a patriot or a traitor.
beatthebrain|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
theknottybride|JasonKander|-0.6597|0.213|0.787|0.0|"RT @JasonKander: If we ignore Russian espionage in our election, we embolden other foreign powers to launch similar attacks on every aspect"
Singer77S|smh|-0.5423|0.189|0.811|0.0|Moscow rules? CIA report raises troubling questions about Donald Trump's relationship with Russia  https://t.co/Q828eqW93C via @smh
Singer77S|linkis|-0.5423|0.189|0.811|0.0|Moscow rules? CIA report raises troubling questions about Donald Trump's relationship with Russia  https://t.co/Q828eqW93C via @smh
DeerParkLady|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
NathanFreier|DefenseOne|0.0|0.0|1.0|0.0|RT @DefenseOne: Obama Orders 10-Year Deep Dive into Election Hacking https://t.co/QIH0t8awqU | @DefTechPat https://t.co/66x7iYcz80
NathanFreier|defenseone|0.0|0.0|1.0|0.0|RT @DefenseOne: Obama Orders 10-Year Deep Dive into Election Hacking https://t.co/QIH0t8awqU | @DefTechPat https://t.co/66x7iYcz80
K1er|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
aimee0715|LOLGOP|0.25|0.058|0.846|0.096|RT @LOLGOP: This election is like if A Christmas Carol ended with Scrooge getting a giant tax break paid for by cutting Tiny Tim off Medica
rayyy_charles|Peter_Wehner|0.743|0.0|0.741|0.259|"RT @Peter_Wehner: Rs shrugging off Russian intervention in our election is a perfect illustration of what @JonHaidt refers to as ""motivate"
luissanapacheco|twitter|0.2023|0.0|0.878|0.122|Trump faces first significant post-election pushback from Republicans over CIA report on Russia https://t.co/yM8G1t0eoj
massgamer911|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
razorhead68|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
razorhead68|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
MediaWatchUS1|RepublicanChick|-0.1779|0.082|0.918|0.0|"RT @RepublicanChick: Liberals are accusing Russia of influencing the election. At the same time, liberals enabled citizens of other countri"
StarvingAuthor|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
voilarie85210|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
HalSpencer1|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
molosovsky|ReaderMeter|0.5859|0.0|0.789|0.211|"RT @ReaderMeter: Created a @Wikipedia stub on ""Russian influence on the 2016 United States presidential election. Heres what it looks lik"
s_karmude|AkshayMarathe|-0.8954|0.355|0.6|0.046|"RT @AkshayMarathe: Peak season on in Goa, but no tourists. Locals extremely upset with BJP, want to exact revenge in upcoming election. #de"
Alice16050204|_Makada_|-0.296|0.115|0.826|0.06|"RT @_Makada_: President-Elect Trump: It's ridiculous to say Russia intervened in the election, I think it's just another excuse. We had a m"
ciberjosefina|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
GeorgeHiggins|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
CucusMusic|twitter|0.2023|0.0|0.878|0.122|Trump faces first significant post-election pushback from Republicans over CIA report on Russia https://t.co/lxOpAzgo0Q
ReneeBevevino|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
ReneeBevevino|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
lghcox|Yascha_Mounk|-0.4019|0.119|0.881|0.0|"RT @Yascha_Mounk: German officials: Russia hacked Bundestag, released secret docs, will likely try to influence '17 election as in USA http"
MErb1962|noturbone|0.0|0.0|1.0|0.0|@noturbone https://t.co/uBn6DSJCPt
MErb1962|armed-services|0.0|0.0|1.0|0.0|@noturbone https://t.co/uBn6DSJCPt
AndreFrato|An0nKn0wledge|-0.5859|0.147|0.853|0.0|RT @An0nKn0wledge: They Told Me I Couldn't Have Aliens Hillary &amp; Election Fraud In Same Tweet It Couldn't Be Done They We're Wrong.. http
pgrandee10|IMPL0RABLE|0.0|0.0|1.0|0.0|RT @IMPL0RABLE: #TheResistanceContact @TheJusticeDeptDemand a suppression extension &amp; investigation of election per @CIA concerns of Rus
grt8guy|twitter|-0.7269|0.253|0.747|0.0|Hey Loser even heir Hillary's network said the election could be hacked. #LyingLiberals you cannot have it both way https://t.co/12MdOB2Q5s
ChristineParini|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
ChristineParini|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
dwyer6328|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
KarenCrow6|LeahR77|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
KarenCrow6|t|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
donna980|6bird4|-0.2023|0.116|0.808|0.076|RT @6bird4: @KestrelArts @CaroleDoms @nypost Lost 100% of the presidency. Our forefathers carefully considered our election process https:/
donna980||-0.2023|0.116|0.808|0.076|RT @6bird4: @KestrelArts @CaroleDoms @nypost Lost 100% of the presidency. Our forefathers carefully considered our election process https:/
ji57o|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
KilianJulianus|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/4PzoMvjVdc
Donna_DHKBB|johnastoehr|0.5859|0.0|0.787|0.213|"RT @johnastoehr: FBI covered up Russian influence on Trump's election win, Harry Reid claims https://t.co/UccTvagE8D"
Donna_DHKBB|theguardian|0.5859|0.0|0.787|0.213|"RT @johnastoehr: FBI covered up Russian influence on Trump's election win, Harry Reid claims https://t.co/UccTvagE8D"
clever_monkey|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
mystarisfading|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
SocialCivility|OnlyWhiteTiger|0.0|0.0|1.0|0.0|RT @OnlyWhiteTiger: @JMZElection It should be the entire election including senate and House seats
mindfulzoo|HamiltonElector|0.34|0.0|0.833|0.167|Give CIA Security Briefing to Electors on Russian Election Interference https://t.co/1XXHHktdnd #hamiltonelectors @HamiltonElector
mindfulzoo|petitions|0.34|0.0|0.833|0.167|Give CIA Security Briefing to Electors on Russian Election Interference https://t.co/1XXHHktdnd #hamiltonelectors @HamiltonElector
onthetrail2016|ref|0.0|0.0|1.0|0.0|"SurveyUSA  &amp;raquo; Blog Archive   &amp;raquo; In a Trump vs Clinton Presidential Election, 4 in 10 Voters Will Hold ... https://t.co/onoPiVorSo"
penny63434309|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
therussophile|therussophile|0.5267|0.0|0.673|0.327|Legislature speaker winning presidential election inMoldovas https://t.co/pt1akopJVo https://t.co/yvbOiSVmrd
CJThompson87|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
douglasscraigky|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
douglasscraigky||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
4plaintiff|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
TheOralBuffet|Change|-0.2003|0.121|0.879|0.0|Demand An Audit Of The 2016 Presidential Election - Sign the Petition! https://t.co/cAia02lIPA via @Change
TheOralBuffet|change|-0.2003|0.121|0.879|0.0|Demand An Audit Of The 2016 Presidential Election - Sign the Petition! https://t.co/cAia02lIPA via @Change
deryloconstruct|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
MatthewBParksSr|rwindrem|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
MatthewBParksSr|nbcnews|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
DanielDastti|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
mekmtl|DougHenwood|0.296|0.0|0.804|0.196|RT @DougHenwood: Its ok to manipulate some elections https://t.co/h4ZNsWx1nU https://t.co/HeuenVGwVZ
mekmtl|observer|0.296|0.0|0.804|0.196|RT @DougHenwood: Its ok to manipulate some elections https://t.co/h4ZNsWx1nU https://t.co/HeuenVGwVZ
RubeBait|BruceBartlett|0.0|0.0|1.0|0.0|"RT @BruceBartlett: The question isn't why Russia interfered in our election, the question is why did in interfere on behalf of Trump &amp; the"
ARepublic|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
samiam321123|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
natuphillies|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
TerriLSelby|DailyCaller|-0.3182|0.141|0.859|0.0|RT @DailyCaller: FBI Disagrees With CIA On Russian Influence In The Presidential Election https://t.co/A7trnqgmiA https://t.co/bIIQ5UqyKM
TerriLSelby|dailycaller|-0.3182|0.141|0.859|0.0|RT @DailyCaller: FBI Disagrees With CIA On Russian Influence In The Presidential Election https://t.co/A7trnqgmiA https://t.co/bIIQ5UqyKM
RalphHornsby|youtube|-0.128|0.239|0.541|0.22|Free Speech Under Attack: Deep State Promotes Fake News and False Flag Putin Election Hacking Myths - YouTube https://t.co/JhkYwlSuBv
MarvinKey74|EveningStarNM|0.5413|0.0|0.837|0.163|@EveningStarNM @DarbyKathleen @JoyAnnReid @KTwoSO this election made really inspired me to get involved. this is not over for me
Balthier28|France4Hillary|-0.3612|0.128|0.872|0.0|"RT @France4Hillary: Given @CIA's evidence that Trump rigged the election with Russia, what should happen? #TrumPutingate #RussianHacking #L"
pobandit12|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
bachic2|Amy_Siskind|-0.2023|0.133|0.766|0.101|"RT @Amy_Siskind: It seems like Friday's outrage about the CIA Report and Russia's infiltrating our election, has simmered down to a whimper"
donnaepowell|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
mllnialnews|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
bhaikes|realDonaldTrump|-0.0572|0.058|0.942|0.0|@realDonaldTrump @NBCNightlyNews @CNN So- do you not want to have the briefings b/c they report that Russia interfered with the election?
JenLynnOh|BreitbartNews|-0.822|0.434|0.495|0.071|RT @BreitbartNews: Why do Democrats want a war with Russia so badly? https://t.co/KfMP9vzZsu
JenLynnOh|breitbart|-0.822|0.434|0.495|0.071|RT @BreitbartNews: Why do Democrats want a war with Russia so badly? https://t.co/KfMP9vzZsu
Britneytica|keith_caulfield|0.0|0.0|1.0|0.0|"RT @keith_caulfield: ""McCain, Graham, Schumer, Reed Joint Statement on Reports That Russia Interfered with the 2016 Election"" https://t.co/"
Britneytica|t|0.0|0.0|1.0|0.0|"RT @keith_caulfield: ""McCain, Graham, Schumer, Reed Joint Statement on Reports That Russia Interfered with the 2016 Election"" https://t.co/"
Lwme07|coton_luver|-0.0516|0.162|0.684|0.154|"RT @coton_luver: Supreme Court: Election Can Be Invalidated Due To Massive Fraud, Install Opponent (DETAILS) https://t.co/zIU7YO34mS via @B"
Lwme07|bipartisanreport|-0.0516|0.162|0.684|0.154|"RT @coton_luver: Supreme Court: Election Can Be Invalidated Due To Massive Fraud, Install Opponent (DETAILS) https://t.co/zIU7YO34mS via @B"
DevinKuchynka|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
DevinKuchynka||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
mrsbinker|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
mrsbinker||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
nana2hallie|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
redinfinity|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
redinfinity||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Scribe53|FrankLuntz|-0.3182|0.113|0.887|0.0|RT @FrankLuntz: CIA veterans  none of them fans of Donald Trump  are urging caution about leaked allegations of #RussiaHacking.https:
Coreybez1|dwaynecobb|0.7096|0.0|0.781|0.219|RT @dwaynecobb: ....    So Russia gives election to Trump &amp; Russia gets Tillerson at State and Flynn as National Security Adviser as a bonus
Iam_Books|abuhena0044|-0.1531|0.144|0.693|0.163|RT @abuhena0044: @HamiltonElector _Trump hijacked the election with Russian intervention committing treason to serve multiple interests at
shermsIR|JimGoldgeier|0.2732|0.0|0.909|0.091|"RT @JimGoldgeier: George HW Bush election in '88, the last time Democrats and Republicans alike accepted legitimacy of new POTUS, seems lik"
PennyHunt12|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
RBStalin|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
jannm|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
mtduarte_|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
mtduarte_|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
kingblais|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
ibpixiechick|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
ibpixiechick||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
MissLin68640163|JYSexton|-0.7269|0.268|0.641|0.09|RT @JYSexton: Who cooked intelligence to get a war in Iraq and now have the nerve to go on TV and criticize evidence that Russia hacked our
JoyLightIN|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: @thedailybeast Bernstein also said Comey wouldn't have announced pre-election unless something major. Woodward said ema
AdrianF1erros|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
SarahsMimi|quinncy|-0.25|0.136|0.777|0.087|RT @quinncy: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/98YVepksgE via @PalmerR
SarahsMimi|palmerreport|-0.25|0.136|0.777|0.087|RT @quinncy: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/98YVepksgE via @PalmerR
Teelin|DarkoftheWeb|0.3612|0.0|0.815|0.185|@DarkoftheWeb *at the end of the yarn is an election cycle* :-p
DannettaJohnson|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
azpat0|youtube|-0.7865|0.409|0.591|0.0|CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia https://t.co/048RfmUA1E
dr_bruin|bros4hillary|0.0|0.0|1.0|0.0|Daily Digest - Election Watch 2016 https://t.co/kDjOfv6DMI via @bros4hillary
dr_bruin|linkis|0.0|0.0|1.0|0.0|Daily Digest - Election Watch 2016 https://t.co/kDjOfv6DMI via @bros4hillary
anobscureartist|casatino|-0.1027|0.097|0.903|0.0|RT @casatino: FBI: sends vague letter; actually nothingMSM: *quivers*CIA: confirms Russia interfered w/electionMSM: \_()_/https://
ryanhide|zandywithaz|-0.3182|0.095|0.905|0.0|@zandywithaz If the election were held 2 weeks earlier she probably just loses a chunk of her pop vote lead. He had a ROUGH last 2 weeks.
macmcd|HRCNJVolunteers|0.3164|0.0|0.887|0.113|RT @HRCNJVolunteers: @GoddessKerriLyn Little sense in 2nd election while Russia's hacking. &amp; another chance to vote for Russia Colluder?! N
AgQueue|armed-services|0.0|0.0|1.0|0.0|"McCain, Graham, Schumer, Reed Joint Statement on Reports That Russia Interfered with 2016 Election https://t.co/QU4rUK8aTI"
teqminsky|change|0.4215|0.0|0.865|0.135|"In light of recent evidence reported by the CIA, that the United States 2016 Presidential Election has been... https://t.co/leIe39klc1"
ElenaSryva|eileendefreest|0.0|0.0|1.0|0.0|"RT @eileendefreest: #ImStillNotOver the fact that Trump, Comey, and GOP Congress aren't in jail yet for allowing Russia to decide the elect"
sstuart2016|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
sstuart2016|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
fuddrucker1|jabeale|0.4019|0.0|0.881|0.119|"RT @jabeale: If Russia clandestinely interfered with a US election in order to favor a particular candidate, POTUS and the CIA should make"
mswindy12|Shoq|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
mswindy12|t|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
PatDugan|LeahR77|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
PatDugan|t|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
AbsP|sacca|0.6369|0.088|0.654|0.258|RT @sacca: On @NPR I shared why tech leaders who go to Trump Tower will get played and also lose the respect of employees. https://t.co/XGA
AbsP|t|0.6369|0.088|0.654|0.258|RT @sacca: On @NPR I shared why tech leaders who go to Trump Tower will get played and also lose the respect of employees. https://t.co/XGA
deleonora_abel|GeorgeTakei|0.34|0.0|0.902|0.098|"RT @GeorgeTakei: If there was interference on the play, you don't count the touchdown. Russia meddled in our election, says the CIA. Electo"
iveygirl08|topbuzzapp|0.0|0.0|1.0|0.0|Latest Election Results: Congressman Calls On Elec... https://t.co/ogI6BIHWxp
DeerParkLady|TrumpsNewsDaily|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
DeerParkLady|yahoo|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
weezmgk|robreiner|0.0|0.0|1.0|0.0|"RT @robreiner: Teapot Dome,Watergate,Iran-Contra are quaint compared to Russian gov. in league with Trump to influence US election. Crimina"
Roxy4080|SpyTalker|0.4767|0.0|0.795|0.205|RT @SpyTalker: CIA Veterans Urge Immediate all-agency National Intelligence Estimate on Trump-Russia https://t.co/Wv2ZCpd0Yw
Roxy4080|newsweek|0.4767|0.0|0.795|0.205|RT @SpyTalker: CIA Veterans Urge Immediate all-agency National Intelligence Estimate on Trump-Russia https://t.co/Wv2ZCpd0Yw
herlipsticklife|leahmcelrath|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
herlipsticklife|t|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
WendiSmith18|slone|0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
WendiSmith18||0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
flgrammardiva|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
scott_stalker2|CarmineZozzora|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
scott_stalker2|t|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
yoshinofarmky|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
yoshinofarmky|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
jmood88|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
urbanista01|Valeriegromes16|0.6351|0.0|0.827|0.173|"@Valeriegromes16 Hahaha, what are you even talking about?! You're cracking me up! The election is over. Now it's about putting #AmericaFirst"
Mellecon|noisyparker|-0.631|0.179|0.821|0.0|"RT @noisyparker: @Mellecon Youd think theyd be extra-sensitive about that post-election, but it never enters their head that ""fake news"
mowser1970|foxnation|0.0|0.0|1.0|0.0|"RT @foxnation: .@JudgeJeanine: The Election Is Over, Mr. President https://t.co/VW0vBabMjz"
mowser1970|nation|0.0|0.0|1.0|0.0|"RT @foxnation: .@JudgeJeanine: The Election Is Over, Mr. President https://t.co/VW0vBabMjz"
vinyldude82|_Makada_|0.0431|0.113|0.768|0.119|"RT @_Makada_: Obama ordered intelligence agencies to investigate Russian interference in election with NO PROOF, by doing this he is the on"
Cnvido|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
rosereynolds|NoceraNYT|0.0|0.0|1.0|0.0|RT @NoceraNYT: Is this for real?  https://t.co/AHODO2pTpa
rosereynolds|palmerreport|0.0|0.0|1.0|0.0|RT @NoceraNYT: Is this for real?  https://t.co/AHODO2pTpa
Rink_Mama|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
ActorAaronBooth|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
m364np4163|ParkerMolloy|-0.5067|0.17|0.83|0.0|"RT @ParkerMolloy: ""patrioteagle.flag says there's a child sex pizza dungeon!""""On it!""""The CIA says Russia messed w/ the election!""Some s"
jtvrdik|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
PennyFate|twitter|-0.296|0.141|0.763|0.095|7/we can have fruit from the poisonous tree. One remark to you. This election has bent the rules like never before. https://t.co/wglTb65sTk
ohaginib|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ToddFleming123|LindaSuhler|-0.2168|0.144|0.75|0.106|RT @LindaSuhler: Remember Obama's hot mic msg to Putin about flexibility after the election?What are they scared of? #RussianHackinghttps
Gregorylund|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
sarefo|leahmcelrath|0.5584|0.0|0.796|0.204|RT @leahmcelrath: Watergate seems like such an minor almost innocent bit of subterfuge compared to what's happened in this election.
Eonkidz|RealAlexJones|-0.7865|0.348|0.652|0.0|RT @RealAlexJones: #CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia - https://t.co/eXe3mPaIEG #infowars
Eonkidz|youtube|-0.7865|0.348|0.652|0.0|RT @RealAlexJones: #CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia - https://t.co/eXe3mPaIEG #infowars
Peacepox|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
ShencoRR|neil1pat|-0.5859|0.213|0.787|0.0|"RT @neil1pat: Where Tory election fraud claims are being investigated, in one map https://t.co/JkNITwT57b #toryelectionfraud"
ShencoRR|indy100|-0.5859|0.213|0.787|0.0|"RT @neil1pat: Where Tory election fraud claims are being investigated, in one map https://t.co/JkNITwT57b #toryelectionfraud"
StewrtSmthRadio|gourmetspud|-0.7717|0.3|0.7|0.0|"RT @gourmetspud: ""Hillary lost bc fake news"" seems 100x less plausible than ""Hillary lost because she was Democratic Romney in anger-driven"
ChicagoMGD|jkarsh|0.4576|0.0|0.87|0.13|"RT @jkarsh: Given the CIA report about Russia influencing our election, this line from an @azcentral piece is very interesting. https://t.c"
ChicagoMGD||0.4576|0.0|0.87|0.13|"RT @jkarsh: Given the CIA report about Russia influencing our election, this line from an @azcentral piece is very interesting. https://t.c"
Plumazul|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
Plumazul||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
saygnitegracie3|kerrywashington|0.0|0.0|1.0|0.0|@kerrywashington Total Recount and Audit! Chuck Schumer calls for probe into Russian interference in the election
Alllwftopic|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
erin_d9|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
BevPerryMusic|nytimes|-0.7096|0.258|0.742|0.0|RT @nytimes: Donald Trump ties CIA reports on Russian meddling in the election to Democrats' embarrassment over defeat https://t.co/2QMNlJ3
BevPerryMusic|t|-0.7096|0.258|0.742|0.0|RT @nytimes: Donald Trump ties CIA reports on Russian meddling in the election to Democrats' embarrassment over defeat https://t.co/2QMNlJ3
BourneInTexas|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
Marypat714|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
Rink_Mama|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
L188188|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
BamaStephen|DavidAFrench|-0.3612|0.122|0.878|0.0|RT @DavidAFrench: What's the argument against a bipartisan investigation of Russian efforts to disrupt and/or influence the election? Is th
TeamTrumpTeX|ShennaFoxMusic|0.0772|0.0|0.929|0.071|"RT @ShennaFoxMusic: Russia intervened in election #PresidentElect ""Ridiculous, just another excuse, Dems pushing the story, WE had a massiv"
nopocketspapi|ratcake655321|-0.3182|0.084|0.916|0.0|"@ratcake655321 in a nutshell, if you such a lack of use for an ID that you don't have one, the effect of the election on you is negligible."
art_f2001|Allnkat|-0.2732|0.126|0.754|0.121|RT @Allnkat: She is laughable:         Kellyanne Conway calls CIA report on Russian election meddling laughable and ridiculous https://t.
art_f2001||-0.2732|0.126|0.754|0.121|RT @Allnkat: She is laughable:         Kellyanne Conway calls CIA report on Russian election meddling laughable and ridiculous https://t.
aplemkseriously|BruceBartlett|0.0|0.0|1.0|0.0|"RT @BruceBartlett: The question isn't why Russia interfered in our election, the question is why did in interfere on behalf of Trump &amp; the"
surfsalterpath|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
surfsalterpath|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
greggwall|twitter|0.7259|0.0|0.783|0.217|Election is old news. Obama is old news. Pres Elect Trump only wants what is best for us not worried about old news https://t.co/rZdAKpwocY
kysgabbygirl|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
ClintCastleford|nationalpost|-0.3612|0.161|0.839|0.0|Donald Trump says its ridiculous to think Russia interfered in election https://t.co/nHPUpUtsEk via @nationalpost
ClintCastleford|news|-0.3612|0.161|0.839|0.0|Donald Trump says its ridiculous to think Russia interfered in election https://t.co/nHPUpUtsEk via @nationalpost
PolitixGal|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
PolitixGal|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
mgyousey|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
mgyousey|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
shaqueelsinai|ianbremmer|-0.34|0.107|0.893|0.0|RT @ianbremmer: I don't believe Russia intervention changed the outcome of election. But to deny CIA evidence of direct hacking is traito
rhenderson7110|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
PhilipRWFG|EricBoehlert|0.0|0.0|1.0|0.0|"RT @EricBoehlert: this is why, to date, we have to rely on anonymous sources for information re: Russia and election https://t.co/OSbrbw66M5"
PhilipRWFG|twitter|0.0|0.0|1.0|0.0|"RT @EricBoehlert: this is why, to date, we have to rely on anonymous sources for information re: Russia and election https://t.co/OSbrbw66M5"
Kane_Says405|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
cussetabraswell|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
cussetabraswell||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
_mims16|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
BlackTowerRadio|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
BlackTowerRadio|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
bvkcitizen|KurtSchlichter|-0.1779|0.105|0.817|0.078|RT @KurtSchlichter: You progs can't blow the Russians for four decades then lose an election and convince me you've all of a sudden develop
spzkaz|1Marchella|-0.1531|0.078|0.922|0.0|"RT @1Marchella: ""We've got no evidence that #RussianHackers influenced the election, but we're going to report they did anyway"" https://t.c"
spzkaz||-0.1531|0.078|0.922|0.0|"RT @1Marchella: ""We've got no evidence that #RussianHackers influenced the election, but we're going to report they did anyway"" https://t.c"
TrumpismBook|mathewsjw|-0.6249|0.215|0.785|0.0|RT @mathewsjw: EU Brussels crisis as Le Pen #FranceExit storms into poll lead over rivals  https://t.co/oHzywnokmw
TrumpismBook|express|-0.6249|0.215|0.785|0.0|RT @mathewsjw: EU Brussels crisis as Le Pen #FranceExit storms into poll lead over rivals  https://t.co/oHzywnokmw
bergeronprocess|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
JoanneFralin|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Seacretsoc1|NoceraNYT|0.0|0.0|1.0|0.0|RT @NoceraNYT: Is this for real?  https://t.co/AHODO2pTpa
Seacretsoc1|palmerreport|0.0|0.0|1.0|0.0|RT @NoceraNYT: Is this for real?  https://t.co/AHODO2pTpa
aawestbrook|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
JaguarJake14|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
vrot01|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
lotusbat|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
mplsmike35|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
opelaguila|greenhousenyt|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
opelaguila|t|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
emzorbit|leahmcelrath|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
emzorbit|t|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
maggie805ca|FoxNews|0.0|0.0|1.0|0.0|RT @FoxNews: U.S. markets since election. https://t.co/NRw2LedQ7u
maggie805ca|twitter|0.0|0.0|1.0|0.0|RT @FoxNews: U.S. markets since election. https://t.co/NRw2LedQ7u
SheriHerman10|Counter_info|-0.4019|0.197|0.803|0.0|RT @Counter_info: How To Instantly Tell If Russia Hacked theElection https://t.co/3kwKPyz1RW https://t.co/ZuOftkoUpV
SheriHerman10|counterinformation|-0.4019|0.197|0.803|0.0|RT @Counter_info: How To Instantly Tell If Russia Hacked theElection https://t.co/3kwKPyz1RW https://t.co/ZuOftkoUpV
tellmecandy|Slate|0.5267|0.0|0.793|0.207|RT @Slate: These two shows have been my ideal post-election escapist TV: https://t.co/Iyok2BRWBS https://t.co/ihfKsgmtvG
tellmecandy|slate|0.5267|0.0|0.793|0.207|RT @Slate: These two shows have been my ideal post-election escapist TV: https://t.co/Iyok2BRWBS https://t.co/ihfKsgmtvG
joannanoon|leahmcelrath|0.5584|0.0|0.796|0.204|RT @leahmcelrath: Watergate seems like such an minor almost innocent bit of subterfuge compared to what's happened in this election.
AshgabatCat|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
tomguz|ericgarland|0.7783|0.0|0.736|0.264|RT @ericgarland: And if the winner of a tainted election chooses to stand against national interest and for that foreign aggressor:The wo
SFDoug|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
amandablount2|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
Apipwhisperer|ShennaFoxMusic|0.0772|0.0|0.929|0.071|"RT @ShennaFoxMusic: Russia intervened in election #PresidentElect ""Ridiculous, just another excuse, Dems pushing the story, WE had a massiv"
coin_seller|ebay|0.0|0.0|1.0|0.0| 1972 McGOVERY EAGLETON 1 1/2 INCH PRESIDENTIAL ELECTION  BUTTON P159 https://t.co/CwUHPoHk7Q https://t.co/yuMS6KxOGk
KelleyEltzroth|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
KelleyEltzroth||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Jasavage76Joyce|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
Jasavage76Joyce||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
mowser1970|FoxNews|0.1027|0.089|0.806|0.105|"RT @FoxNews: Last night on ""Justice,"" @JudgeJeanine had stark words for those who refuse to accept the results of the election. https://t.c"
mowser1970||0.1027|0.089|0.806|0.105|"RT @FoxNews: Last night on ""Justice,"" @JudgeJeanine had stark words for those who refuse to accept the results of the election. https://t.c"
ydavey|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
OakCliffITGuy|NicholsUprising|0.0|0.0|1.0|0.0|"RT @NicholsUprising: ""I believe electors have the right to consider that.""-- US Rep. David Cicilline, D-RI, on potential hacking of electi"
oopsycharlie|JoyceDiDonato|-0.4019|0.206|0.67|0.124|"@JoyceDiDonato Which composer and singers, dead or alive, would you choose for Election 2016: The Opera?"
ActorAaronBooth|GeorgeTakei|-0.4199|0.108|0.892|0.0|"RT @GeorgeTakei: Mitch McConnell tried to cast doubt on the CIA findings before the election. Then, magic! His wife Elaine Chao is named Tr"
gustergrl03|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
charlescollier|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
What_you_sow|Bill_Rhodes54|-0.5994|0.253|0.653|0.094|RT @Bill_Rhodes54: Dems: Russia hacked the electionPatriot: Really how so?Dems: They told Americans the Truth about our horrible candid
KathrynECramer|jacklgoldsmith|0.6124|0.0|0.75|0.25|"RT @jacklgoldsmith: Outstanding, sober account of latest goings-on w Russia and US election.   https://t.co/dtx6Suetfg"
KathrynECramer|nytimes|0.6124|0.0|0.75|0.25|"RT @jacklgoldsmith: Outstanding, sober account of latest goings-on w Russia and US election.   https://t.co/dtx6Suetfg"
FieryRedReviews|twitter|0.0|0.0|1.0|0.0|"The executive branch has called for investigation, and at least one Congressman is calling for a new election. https://t.co/T5LW2dSPV1"
RagingBull300|greenhousenyt|-0.0516|0.11|0.787|0.102|"RT @greenhousenyt: ""The fact that 59% of the vote-counting machines in Detroit all broke on Nov. 8 stands out as a stunning developmnt"" htt"
SeanCollinsCali|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ngelKisses|Reuters|0.0|0.0|1.0|0.0|RT @Reuters: Trump says reports Russia helped him in U.S. election are 'ridiculous' https://t.co/rXNYe3xLYB https://t.co/KahIv6TwG7
ngelKisses|reuters|0.0|0.0|1.0|0.0|RT @Reuters: Trump says reports Russia helped him in U.S. election are 'ridiculous' https://t.co/rXNYe3xLYB https://t.co/KahIv6TwG7
ibpixiechick|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
ibpixiechick|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
Deanna_MG|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
donailin|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
donailin|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Zenkitty714|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
siddharthainc|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
siddharthainc|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
BelisaDavis|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
Jackanaples|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
onlyonebran|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
onlyonebran|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
hyperlocavore|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
iamrami1996|CNN|-0.5106|0.18|0.82|0.0|RT @CNN: Where's the outrage over Russia's hack of the US election? -via @CNNOpinion https://t.co/Rs4QzciIQS https://t.co/DPQ2QJZZVe
iamrami1996|cnn|-0.5106|0.18|0.82|0.0|RT @CNN: Where's the outrage over Russia's hack of the US election? -via @CNNOpinion https://t.co/Rs4QzciIQS https://t.co/DPQ2QJZZVe
carlckitchen|MichaelBKelley|0.0|0.0|1.0|0.0|RT @MichaelBKelley: WikiLeaks seems to be conflating itself with Russian hacking here. Story doesn't mention WikiLeaks. Mask slippage? http
PeabsLord|mattmfm|-0.25|0.274|0.516|0.21|RT @mattmfm: Kellyanne Conway is such a bitter loser. Makes sense when:- you massively lost popular vote- Comey won you election- Russia
andyfroemke1|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
sexxymama131970|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
languageNhumor|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
Clio_On_Kinja|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
VinnieVinnieo|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
JaneMoss08|JuddLegum|0.4404|0.0|0.847|0.153|RT @JuddLegum: Updated list of GOP members supporting investigation into Russian interference w/prez electionSen GrahamSen McCainSen Co
Michael26222747|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
jmerrick82yaho1|twitter|-0.7003|0.327|0.673|0.0|Irony of complaints about foreign involvement in election after the deception of foundation money laundering. Compl https://t.co/5ERWjrEiId
ZeroUtopia|PattyMurray|0.3182|0.0|0.905|0.095|RT @PattyMurray: An investigation must begin as soon as possible on any evidence Russia actively worked to hijack our election &amp; elect Dona
LisaMendoza63|HawaiiDelilah|0.4023|0.0|0.875|0.125|"RT @HawaiiDelilah: Re: Russian interference into our election.If this clip does not outrage you, then you're not paying attention:  https"
to_suesmall|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
aplemkseriously|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
erinpeloso|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
erinpeloso||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
NicoleOrosco4|An0nKn0wledge|-0.5859|0.147|0.853|0.0|RT @An0nKn0wledge: They Told Me I Couldn't Have Aliens Hillary &amp; Election Fraud In Same Tweet It Couldn't Be Done They We're Wrong.. http
AmericanLizzy|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
bonniemac52|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
mariebayarea4|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: @thedailybeast Bernstein also said Comey wouldn't have announced pre-election unless something major. Woodward said ema
tcynthe|SandraRose)I'm|0.0|0.0|1.0|0.0|Retweeted Sandra Rose (@SandraRose):I'm guessing that the majority of Obama's 2008 election campaign donations... https://t.co/GHt5KK7tZY
tcynthe|facebook|0.0|0.0|1.0|0.0|Retweeted Sandra Rose (@SandraRose):I'm guessing that the majority of Obama's 2008 election campaign donations... https://t.co/GHt5KK7tZY
2000Thb|louloubabba|0.5859|0.0|0.787|0.213|"@louloubabba @YouTube Wow, qu'elle pense profonde. L'lection de Trump, un lment du retour des nations"
_coleoptera_|AliMaadelat|0.0|0.0|1.0|0.0|"RT @AliMaadelat: Election People: ""Mr. Trump, you did it! You're going to be President!""Trump: ""Oh... no..."" https://t.co/RQLRJ42KaM"
_coleoptera_|twitter|0.0|0.0|1.0|0.0|"RT @AliMaadelat: Election People: ""Mr. Trump, you did it! You're going to be President!""Trump: ""Oh... no..."" https://t.co/RQLRJ42KaM"
valeyrie47|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
valeyrie47|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
ZeroShits2Give|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
TimerUsa|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
saintwalker98|PattyMurray|0.3182|0.0|0.905|0.095|RT @PattyMurray: An investigation must begin as soon as possible on any evidence Russia actively worked to hijack our election &amp; elect Dona
GENIOCRATIC|bretterlich|-0.5267|0.159|0.841|0.0|.@bretterlich @johniadarola do you realize that it's CENK who is pushing the conspiracy theory that Russia controlled electionNot AlexJones
Allwaysrite55|GartrellLinda|-0.4588|0.136|0.864|0.0|RT @GartrellLinda: Where was @SenJohnMcCain speaking up when obama used taxpayer $ to defeat PM Netanyahu? obama interfered in Israeli elec
artspeaks_|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
artspeaks_||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
DBR96A|d_fucile|-0.5449|0.133|0.867|0.0|RT @d_fucile: THERE'S NO NEW ELECTION!  THE RUSSIANS DIDN'T HACK! ONE MAN WHO WAS INVOLVED WITH ASSANGE ALREADY SAID IT WAS NOT RUSSIANS AS
Ruthperricone|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
TheMrsDarcy|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
AylorKim|FitzyGFY|-0.7574|0.319|0.681|0.0|RT @FitzyGFY: I'm w/@mtdisme - Russia absolutely hacked into Steelers PSI last week to distract from US election accusations #DeflateGate2
ARepublic|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
ARepublic|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
Deemoney521|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
Deemoney521|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
malakim2099|PattyMurray|0.3182|0.0|0.905|0.095|RT @PattyMurray: An investigation must begin as soon as possible on any evidence Russia actively worked to hijack our election &amp; elect Dona
dayy_jay|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
silverkingg|cctvnews|-0.3612|0.135|0.865|0.0|RT @cctvnews: Donald Trump: CIA assessment of Russian interference in US election ridiculous. Follow us for updates.
58isthenew40|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
AkaMotherto3|twitter|-0.4588|0.231|0.769|0.0|Further proof Russia interfered in election. Theyre attacking all democracies. https://t.co/qmtscpG435
tcynthe|SandraRose|0.0|0.0|1.0|0.0|RT @SandraRose: I'm guessing that the majority of Obama's 2008 election campaign donations coming from Saudi Arabia had nothing to do with
michaels_leigh|JamesComeyFBI|-0.2671|0.261|0.568|0.171|Not only does @JamesComeyFBI need to resign We NEED a NEW Election...this one Really Sucked! THANKS 2 https://t.co/FdL5xwDD5S
michaels_leigh|twitter|-0.2671|0.261|0.568|0.171|Not only does @JamesComeyFBI need to resign We NEED a NEW Election...this one Really Sucked! THANKS 2 https://t.co/FdL5xwDD5S
chanale16|BruceBartlett|0.0|0.0|1.0|0.0|"RT @BruceBartlett: The question isn't why Russia interfered in our election, the question is why did in interfere on behalf of Trump &amp; the"
vincedorsett1|thehill|0.0|0.0|1.0|0.0|FBI breaks with CIA on Russia interference in U.S. election https://t.co/AitDIO6DQD
SashaFierce60|MMFlint|0.8689|0.077|0.568|0.355|RT @MMFlint: The CIA has determined Russia hacked into our election to help elect Donald J. Trump. Now Trump names Putin best friend as OUR
bryoneill11|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
djustice7|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
PatDugan|laurahollis61|-0.6486|0.238|0.762|0.0|"RT @laurahollis61: This whole ""Russians hacked the election"" story is the biggest load of crap since#Benghazi ""it-was-a-video."" Dems are d"
thegaf|PattyMurray|0.3182|0.0|0.905|0.095|RT @PattyMurray: An investigation must begin as soon as possible on any evidence Russia actively worked to hijack our election &amp; elect Dona
Noah_Weisberg|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Noah_Weisberg||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
gailmkru|greenhousenyt|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
gailmkru|t|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
ejgabriel9|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
awexton|ndrew_lawrence|-0.128|0.094|0.833|0.072|RT @ndrew_lawrence: Just making sure I've got this rightStarbucks cups and cereal are a reason for outrage but foreign interference in ou
Zoraida12098036|DailyNewsBin|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
Zoraida12098036|palmerreport|-0.3612|0.135|0.865|0.0|"RT @DailyNewsBin: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/LCAfgvCGeY"
EDee_1|JBurtonXP|-0.4019|0.124|0.876|0.0|"RT @JBurtonXP: Always remember that by ""hacked the election,"" these people mean ""released 100% authentic documents that showed real Democra"
devincomiskey|michaelianblack|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
devincomiskey|twitter|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
MobiLibrarian|LibraryJournal|-0.5719|0.198|0.802|0.0|RT @LibraryJournal: New Reference Database: Hate Index: Tracking the Toll of Intolerance Post-Election 2016 https://t.co/Fr9dTTazeR https
MobiLibrarian|infodocket|-0.5719|0.198|0.802|0.0|RT @LibraryJournal: New Reference Database: Hate Index: Tracking the Toll of Intolerance Post-Election 2016 https://t.co/Fr9dTTazeR https
JBax52|theonlyadult|-0.3164|0.098|0.902|0.0|RT @theonlyadult: The noise you just heard is the popping of a vein in my forehead. Cancel the fucking election results now! https://t.co/8
JBax52|twitter|-0.3164|0.098|0.902|0.0|RT @theonlyadult: The noise you just heard is the popping of a vein in my forehead. Cancel the fucking election results now! https://t.co/8
realheine|An0nKn0wledge|-0.6908|0.289|0.619|0.093|RT @An0nKn0wledge: Crazy Thought What If The CIA Yelled #RussiaHacking To Distract From REAL Election Fraud In Favor Hillary &amp; DHS Attempte
sammelbis1998|Kira_G_O_T_N_W|-0.7003|0.358|0.55|0.092|RT @Kira_G_O_T_N_W: Shock poll predicts French Socialists have no chance of beating Marine Le Pen https://t.co/dvExK0kAIV
sammelbis1998|express|-0.7003|0.358|0.55|0.092|RT @Kira_G_O_T_N_W: Shock poll predicts French Socialists have no chance of beating Marine Le Pen https://t.co/dvExK0kAIV
Tracy_Mack|WalshFreedom|0.3182|0.0|0.897|0.103|RT @WalshFreedom: It's not about re litigating the election. It's about finding out what happened. Making sure it never happens againWe s
kwtmobilesalon|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Ronda524|MtnMD|0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
Ronda524||0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
Raj_Bisht5|Dev_Fadnavis|0.0|0.0|1.0|0.0|"RT @Dev_Fadnavis: You voted us in VidhaSabha election;we gave Minister from Nilanga.Now,its time to again vote for #BJP &amp;electNagaradhyaks"
Breruizg|nytimesworld|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
Breruizg|nytimes|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
saadmohseni|ianbremmer|-0.34|0.107|0.893|0.0|RT @ianbremmer: I don't believe Russia intervention changed the outcome of election. But to deny CIA evidence of direct hacking is traito
klormpster|RealAlexJones|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
klormpster|infowars|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
ColinMacKeen|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
classygal21|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
cu_mr2ducks|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
cu_mr2ducks|t|0.0|0.0|1.0|0.0|RT @wikileaks: What was on people's minds about Hillary Clinton during the lead up to the US election? (interactive graph) https://t.co/ts8
Skwidj|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
Skwidj|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
sparkyNadine|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
DarfishIzady|TrumpGo_2016|-0.3182|0.141|0.859|0.0|RT @TrumpGo_2016: FBI Disagrees With CIA On Russian Influence In The Presidential Election https://t.co/nhQAIdZjDX https://t.co/q80zSiwCzZ
DarfishIzady|dailycaller|-0.3182|0.141|0.859|0.0|RT @TrumpGo_2016: FBI Disagrees With CIA On Russian Influence In The Presidential Election https://t.co/nhQAIdZjDX https://t.co/q80zSiwCzZ
Murphy133|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
HillaryWonFools|NewDay|-0.3612|0.161|0.839|0.0|@NewDay you're just further making the case that the election was rigged by Russia....
steelyweather|leahmcelrath|0.5584|0.0|0.796|0.204|RT @leahmcelrath: Watergate seems like such an minor almost innocent bit of subterfuge compared to what's happened in this election.
tkcoffey77|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
genuke1|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
mentalfracking|PalmerReport|-0.7798|0.326|0.598|0.077|Michigan officials admit majority of WTF! Detroit #vote counting machines broke on #Election Day https://t.co/54O22Ff8mb via @PalmerReport
mentalfracking|palmerreport|-0.7798|0.326|0.598|0.077|Michigan officials admit majority of WTF! Detroit #vote counting machines broke on #Election Day https://t.co/54O22Ff8mb via @PalmerReport
fuklikeme|EscapeVelo|-0.3182|0.113|0.887|0.0|RT @EscapeVelo: The FBI leaked that #GamerGate was a Russian psyops operation designed to influence the 2016 Presidential Election. #Stop
LRD90|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Tainoman55|palmerreport|-0.25|0.151|0.753|0.097|Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/64v9bBXYWp via PalmerReport
e_revolutionist|kflana|0.0772|0.116|0.756|0.129|RT @kflana: when you're having a good time and you suddenly remember that you're still upset about the election https://t.co/2GO8TzgJiP
e_revolutionist|twitter|0.0772|0.116|0.756|0.129|RT @kflana: when you're having a good time and you suddenly remember that you're still upset about the election https://t.co/2GO8TzgJiP
ejbshaw|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
lkdavolos|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
lkdavolos||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
otaconred88|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Ericdombro|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
mar82347254|JuddLegum|0.4404|0.0|0.847|0.153|RT @JuddLegum: Updated list of GOP members supporting investigation into Russian interference w/prez electionSen GrahamSen McCainSen Co
wtf_imtooold|Green_Footballs|0.25|0.1|0.72|0.18|RT @Green_Footballs: One thing was confirmed beyond any doubt in this election: the Republican Party is just fine with white supremacism.
Rawkuz99|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
mmmm1026|Khanoisseur|-0.2263|0.087|0.913|0.0|RT @Khanoisseur: More new evidence that Comey tipped undecided voters toward Trump in last 2 weeks of the electionBiggest tamperer was th
B_H_Fan4Evr|IAMKPSmith|0.0|0.0|1.0|0.0|RT @IAMKPSmith: I remember election night kept saying it's all going to come down to Michigan. This is something right out of #scandal.
maxthegirl|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
ginanotjenna|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
theDailyGlobals|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/YAV3H4NGpJ
netminnow|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
pinkbiscuit|MartinWiener|0.0|0.0|1.0|0.0|"RT @MartinWiener: @DENVERSMKC @VictorB123 @brassmonkey3434 If there was proof Obama would have been all over it then, not five weeks after"
gabey8|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
gabey8||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
sluttycatlady|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
FailuresArt|kurteichenwald|0.7906|0.0|0.704|0.296|@kurteichenwald Thank you for your excellent work covering the biggest story of the year about Russian efforts in the US election. Important
PaulMick|ACNewman|0.34|0.124|0.659|0.217|"RT @ACNewman: Look, more shadiness in the election. If true, Michigan was stolen. If that's true, why not others ? https://t.co/OSorsOpmO0"
PaulMick|palmerreport|0.34|0.124|0.659|0.217|"RT @ACNewman: Look, more shadiness in the election. If true, Michigan was stolen. If that's true, why not others ? https://t.co/OSorsOpmO0"
darren_nicholls|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
wmarianne77|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
pjmcgovern4|owillis|-0.296|0.115|0.885|0.0|"RT @owillis: shorter @realDonaldTrump ""if i tweet this maybe thell stop talking about putin buying me an election"" https://t.co/nNttUQHea6"
pjmcgovern4|oliverwillis|-0.296|0.115|0.885|0.0|"RT @owillis: shorter @realDonaldTrump ""if i tweet this maybe thell stop talking about putin buying me an election"" https://t.co/nNttUQHea6"
macmcd|webcodepro|-0.1655|0.145|0.698|0.157|"RT @webcodepro: @GoddessKerriLyn I'd love this to be true, but fake news happens on both sides, will wait &amp; see. There's a Petition https:/"
macmcd||-0.1655|0.145|0.698|0.157|"RT @webcodepro: @GoddessKerriLyn I'd love this to be true, but fake news happens on both sides, will wait &amp; see. There's a Petition https:/"
ashmalaviya|nytimes|0.3182|0.0|0.905|0.095|This explains the election results in the USA :-) -&gt; High on Hitler and Meth: Book Says Nazis Were Fueled by Drugs https://t.co/DIpq334KXm
JayDotson__|mikeyymike78|0.0|0.0|1.0|0.0|RT @mikeyymike78: Major week in American politics coming up: Sec of State to be announced amid furor over reports Russia attempted to aide
zone_202|lordaedonis|0.0|0.0|1.0|0.0|RT @lordaedonis: I wonder what it was about the 2016 election that made the russians decide to finally activate 'Operation Make America Gre
JiriLeniValenta|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
CoreyPeper|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
CoreyPeper|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
oscarfc0311|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
SamScrogg|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
BombsTruth|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
Roxy4080|MalcolmNance|0.1027|0.113|0.756|0.13|RT @MalcolmNance: READ: My Spy Thriller-paced book. How Russian Intelligence Hacked the 2016 Election to elect Donald Trump President. http
BananaHeadLady|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
BananaHeadLady||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Katherine022610|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
saksivas_|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
DHeber|nytimes|0.4939|0.0|0.61|0.39|Russias Hand in Americas Election https://t.co/mYfwRlsbkb
AngelinaSnow007|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
NYtitanic1999|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
NYtitanic1999|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
sammelbis1998|mathewsjw|-0.6249|0.215|0.785|0.0|RT @mathewsjw: EU Brussels crisis as Le Pen #FranceExit storms into poll lead over rivals  https://t.co/oHzywnokmw
sammelbis1998|express|-0.6249|0.215|0.785|0.0|RT @mathewsjw: EU Brussels crisis as Le Pen #FranceExit storms into poll lead over rivals  https://t.co/oHzywnokmw
BettinaAnter|greenhousenyt|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
BettinaAnter|t|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
szipster|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
TilloTill|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
darrintyler29|BardockObama|-0.8208|0.322|0.591|0.087|"RT @BardockObama: Liberals are so stupid y'all ask for a recount then fail, then think Russia rigged the election lol it was obviously J Co"
Iamnowblue|emigre80|-0.3802|0.217|0.662|0.121|"RT @emigre80: Both Trump and Sanders were delighted to cry ""rigged election!"" when they ran against Clinton.Now that there's evidence? *C"
CreativeArtAPE|freddiedeboer|0.34|0.0|0.888|0.112|"RT @freddiedeboer: The most striking, consistent aspect of post-election behavior from Democrats is the absolute refusal to engage in real"
JeffCallahan75|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
JeffCallahan75|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
slickvolt|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
slickvolt|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
MichaelTetrick|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
kwtmobilesalon|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
ggnewsus|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/DhMMngCm1J
Atticus_Amber|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
marcel_g|sproudfoot|0.0|0.0|1.0|0.0|"RT @sproudfoot: This is an absolute tour de force. On game theory, Russia and the election: https://t.co/o6LOUq36P9"
marcel_g|storify|0.0|0.0|1.0|0.0|"RT @sproudfoot: This is an absolute tour de force. On game theory, Russia and the election: https://t.co/o6LOUq36P9"
pdevhecht|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
pdevhecht|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
rogiloc|DatPissedOffCat|-0.296|0.136|0.864|0.0|RT @DatPissedOffCat: @LindseyGrahamSC @SenSchumer @SenJohnMcCain This was an #InvalidElection #RevoteNow No #inauguration for ANYONE till t
e_revolutionist|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
richeagle100|BreitbartNews|-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
richeagle100||-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
randalltrandall|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
Vinogamist|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
Vinogamist|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
devanieangel|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
jvargasnow|TroyBlayne|-0.3182|0.139|0.772|0.089|RT @TroyBlayne: @guypbenson @jvargasnow @Zegota42 It would be illegal for the CIA to be actively working to interfere or disrupt the electi
maderaedwards|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
lolaa1956|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
benhaygood|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
AliciaGs_BigMa|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
Betterw05759703|AtticusinCanada|0.0|0.0|1.0|0.0|RT @AtticusinCanada: @amjoyshow @debilu2 @SenatorReid He absolutely should be. They gamed the election on purpose using Comey.
rdsono|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
JHowieJr|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
JwchrisJon|jaketapper|-0.4404|0.178|0.822|0.0|@jaketapper Delay Trump taking office until it can be verified to what extent the hacking affected the election. Remember 2000
Spacekatgal|PattyMurray|0.3182|0.0|0.905|0.095|RT @PattyMurray: An investigation must begin as soon as possible on any evidence Russia actively worked to hijack our election &amp; elect Dona
INVUQT|cristinalaila1|0.0|0.0|1.0|0.0|RT @cristinalaila1: MSM is more concerned about unsubstantiated claims of Russia hacking the election than Hillary's maid printing up class
ikengachronicle|twitter|0.0|0.0|1.0|0.0|Rivers State Election https://t.co/CIuAwhOPcM
LauraK205|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
iblibs|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
mistermichaelk|pixelatedboat|-0.4585|0.167|0.833|0.0|RT @pixelatedboat: I read the 12th Amendment and technically neither Clinton nor Trump won the election: https://t.co/fKieKK3fEH
mistermichaelk|twitter|-0.4585|0.167|0.833|0.0|RT @pixelatedboat: I read the 12th Amendment and technically neither Clinton nor Trump won the election: https://t.co/fKieKK3fEH
JTrachtman|nytimes|0.4939|0.0|0.61|0.39|Russias Hand in Americas Election https://t.co/33noQWNvYf
waltdog4|kurteichenwald|-0.2382|0.22|0.67|0.11|"RT @kurteichenwald: No offense, @chucktodd, but when u say no one was sure Russia behind hack pre-election, shows u need to read more. http"
TeamTrumpTeX|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
207Curtin|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
207Curtin|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
LAKINGSFAN1967|JeffreyGoldberg|0.0534|0.122|0.748|0.129|@JeffreyGoldberg you are a fucking idiot. If there was anything to that story then Obama would have used it during the election for DNC win
tomrichardson80|BrendanNyhan|-0.4659|0.169|0.787|0.043|"RT @BrendanNyhan: Seeing people dismiss as silly conspiracy talk, but far more serious. Potential Dep SOS suggesting Obama used IC in a dom"
gramma61|KeepAmerGr8|-0.5719|0.222|0.778|0.0|RT @KeepAmerGr8: Bipartisan anger grows over Russian interference into U.S. election https://t.co/9MgHpkwma0 via @HuffPostPol
gramma61|huffingtonpost|-0.5719|0.222|0.778|0.0|RT @KeepAmerGr8: Bipartisan anger grows over Russian interference into U.S. election https://t.co/9MgHpkwma0 via @HuffPostPol
jaureguisrivera|danversohara|0.0|0.0|1.0|0.0|RT @danversohara: Everyone around me: the election is over get over itMe: https://t.co/ykfoZyr5k2
jaureguisrivera|twitter|0.0|0.0|1.0|0.0|RT @danversohara: Everyone around me: the election is over get over itMe: https://t.co/ykfoZyr5k2
to_suesmall|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
to_suesmall|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
usa_dmc|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
MissLin68640163|CarisSevern|-0.5719|0.222|0.778|0.0|RT @CarisSevern: Bipartisan anger grows over Russian interference into U.S. election https://t.co/5wkqo8lptj via @HuffPostPol
MissLin68640163|huffingtonpost|-0.5719|0.222|0.778|0.0|RT @CarisSevern: Bipartisan anger grows over Russian interference into U.S. election https://t.co/5wkqo8lptj via @HuffPostPol
FuckJoshura|BardockObama|-0.8208|0.322|0.591|0.087|"RT @BardockObama: Liberals are so stupid y'all ask for a recount then fail, then think Russia rigged the election lol it was obviously J Co"
ambercat7|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
ambercat7|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
simplyhoran|swin24|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
simplyhoran|thedailybeast|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
FishManwaters|FoxNewsSunday|0.0|0.0|1.0|0.0|RT @FoxNewsSunday: Coming up on #FNS -- @realDonaldTrump describes what went through his mind on election night. https://t.co/tJ7myY6Sxk
FishManwaters|twitter|0.0|0.0|1.0|0.0|RT @FoxNewsSunday: Coming up on #FNS -- @realDonaldTrump describes what went through his mind on election night. https://t.co/tJ7myY6Sxk
lawwtey|TrumpsNewsDaily|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
lawwtey|yahoo|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
aplemkseriously|tgreene319|0.0|0.0|1.0|0.0|RT @tgreene319: Let's review. CIA says Russian hackers interfered w election. Russia says they didn't. Trump doesn't believe CIA &amp; instead
bshaurette|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
PaWright10|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
PaWright10|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
jeepeg|europa-news|-0.3612|0.172|0.828|0.0|Donald Trump says CIA charge Russia influenced election is ridiculous | US news https://t.co/5iZ9feHEkV
SharonS72105601|TrumpsNewsDaily|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
SharonS72105601|yahoo|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
lipchikphoto|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
JessicaNexus|mickeybreezy|0.0|0.0|1.0|0.0|@mickeybreezy @Realpolitiki This is my last tweet to you: https://t.co/T6ryyrGejX. You need to read more before the next election.
JessicaNexus|fivethirtyeight|0.0|0.0|1.0|0.0|@mickeybreezy @Realpolitiki This is my last tweet to you: https://t.co/T6ryyrGejX. You need to read more before the next election.
jrussell264|quinncy|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
jrussell264|palmerreport|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
chlotobe|sarahclazarus|0.3182|0.0|0.901|0.099|RT @sarahclazarus: We'll know for sure the Russians were involved if we look into the election and find a smaller election right inside
snarkytoes|VABVOX|0.0|0.0|1.0|0.0|"RT @VABVOX: .@SpeakerRyan is tweeting about overturning #Obamacare, not Russian interference with our election. https://t.co/4SirvxWCKi"
snarkytoes|twitter|0.0|0.0|1.0|0.0|"RT @VABVOX: .@SpeakerRyan is tweeting about overturning #Obamacare, not Russian interference with our election. https://t.co/4SirvxWCKi"
netminnow|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
cussetabraswell|InfoPasser|-0.25|0.136|0.777|0.087|RT @InfoPasser: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/nLL5ZdUfKq via @Palm
cussetabraswell|palmerreport|-0.25|0.136|0.777|0.087|RT @InfoPasser: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/nLL5ZdUfKq via @Palm
blanca10|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
JosephMiller3|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
saksivas_|LeahR77|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
saksivas_|t|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
tom_luu|CNN|0.0|0.0|1.0|0.0|@CNN @inmateschildren 2016 Election Recap: https://t.co/bLhh9FmlTl
tom_luu|twitter|0.0|0.0|1.0|0.0|@CNN @inmateschildren 2016 Election Recap: https://t.co/bLhh9FmlTl
veve4heart|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
susan_424|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
SNetibutr|DebGoBlue|0.0096|0.062|0.875|0.063|RT @DebGoBlue: Once in recess they can't stop it. Well know election secret. Even #bossTrump can't reverse but then #BossTrump is a #fascis
srinivas_vs9|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
formarrowdbs|PatriotGeorgia|-0.5994|0.187|0.813|0.0|RT @PatriotGeorgia: RINO War Hawks Lindsey Graham and John McCain Call for Investigation of Russia Influencing Election https://t.co/EavySu
formarrowdbs|t|-0.5994|0.187|0.813|0.0|RT @PatriotGeorgia: RINO War Hawks Lindsey Graham and John McCain Call for Investigation of Russia Influencing Election https://t.co/EavySu
atgattrat|MaydnUSA|-0.4019|0.119|0.881|0.0|"RT @MaydnUSA: When Sony was hacked, the FBI immediately produced evidence. Anyone seen any actual evidence of election hack by Russia?Did"
povozim|ZimPeopleFirst|-0.6249|0.242|0.758|0.0|@ZimPeopleFirst election agents in Bikita West Struggle Nyahunda &amp; Tsvuru Gurwe beaten up at instigation of Zanu-PF https://t.co/6rk937tHTu
povozim|twitter|-0.6249|0.242|0.758|0.0|@ZimPeopleFirst election agents in Bikita West Struggle Nyahunda &amp; Tsvuru Gurwe beaten up at instigation of Zanu-PF https://t.co/6rk937tHTu
ImCAntonio|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Aszneth|politicususa|-0.7096|0.33|0.67|0.0|Treasonous Mitch McConnell Refused To Oppose Russia Election Meddling For Trump via @politicususa https://t.co/fDXFOHAPIb
Aszneth|politicususa|-0.7096|0.33|0.67|0.0|Treasonous Mitch McConnell Refused To Oppose Russia Election Meddling For Trump via @politicususa https://t.co/fDXFOHAPIb
charles_gaba|MarkBrewerDems|-0.3612|0.102|0.898|0.0|RT @MarkBrewerDems: Time for reform: the legacy of @migop @MichSoS Ruth Johnson is the mess of an election system the recount revealed http
shaylasnali|tgreene319|0.0|0.0|1.0|0.0|RT @tgreene319: Let's review. CIA says Russian hackers interfered w election. Russia says they didn't. Trump doesn't believe CIA &amp; instead
zoegits|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/s1JEK0zXJG
geege4|pattonoswalt|0.4939|0.0|0.882|0.118|"RT @pattonoswalt: Seems to me, you didn't wanna talk about it before the election. Seems to me, you just turned your pretty head &amp; walked a"
Cheerful_7|cerenomri|0.0|0.0|1.0|0.0|"RT @cerenomri: Remember that one week during the election when the left was really, really concerned about anti-Semitism?They're supporti"
OpalescentMoon|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
llh7167|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
llh7167||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
tealalltheway|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
tealalltheway|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
GarthDerby|JasonKander|-0.6597|0.213|0.787|0.0|"RT @JasonKander: If we ignore Russian espionage in our election, we embolden other foreign powers to launch similar attacks on every aspect"
charlesofidaho|ericgarland|0.7783|0.0|0.736|0.264|RT @ericgarland: And if the winner of a tainted election chooses to stand against national interest and for that foreign aggressor:The wo
jonhartmannjazz|t|0.5904|0.0|0.832|0.168|SCOTUS: Invalidate Election Results Of 2016 - Order A New Election https://t.co/zWEJppoFibDO THIS NOW AND GET ALL YOUR FRIENDS TO SIGN NOW
ecstasydragon|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
HH75876116|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
Sgroberts121657|MarieTitus9|-0.1419|0.054|0.946|0.0|@MarieTitus9 I did not agree with his rederick this election but for me and my own we could not or would not go with the same ole same ole
noisyparker|Mellecon|-0.631|0.172|0.828|0.0|"@Mellecon Youd think theyd be extra-sensitive about that post-election, but it never enters their head that ""fake news applies to them."
SentientHunter|GavinNewsom|-0.3089|0.101|0.899|0.0|RT @GavinNewsom: Trump's treating Russian interference in our election as partisan issue. This is not about political parties - our natl se
used2bnew|politico|0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
used2bnew||0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
Lwme07|USARedOrchestra|-0.197|0.098|0.834|0.068|RT @USARedOrchestra: The reason this election didn't seem normal is bcs it wasn't normal so there r no normal solutions. It wasn't an elect
abirish|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
dadavies|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
soldierDtruth|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
JenniferGassman|tgreene319|0.0|0.0|1.0|0.0|RT @tgreene319: Let's review. CIA says Russian hackers interfered w election. Russia says they didn't. Trump doesn't believe CIA &amp; instead
H2E4G|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
H2E4G|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
CALEBHITT|zerohedge|-0.4767|0.162|0.838|0.0|"Joe Scarborough: Hillary Clinton Cost Hillary Clinton the Election, Not Fake News | Zero Hedge https://t.co/5u8ui1TCCq #Trump #Hillary"
MsScree|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
tootropic|Change|0.0|0.0|1.0|0.0|President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/TMSKPRZRsG via @Change
tootropic|change|0.0|0.0|1.0|0.0|President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/TMSKPRZRsG via @Change
TalatAman|sethmoulton|0.6808|0.0|0.811|0.189|"RT @sethmoulton: Proud to see so many #MA6 constituents ready to work for change. There is so much to do, and this election was a call to a"
Sharan116|RealAlexJones|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
Sharan116|infowars|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
hi_hat_truth|neeratanden|0.0|0.0|1.0|0.0|@neeratanden @EricLiptonNYT @ScottShaneNYT @EricLichtblau @nytimes why are the election results still being considered valid?
simplyhoran|swin24|-0.0572|0.055|0.945|0.0|"RT @swin24: Today, Trump says he doesnt want anyone hacking the U.S.In July, he called on Russia to hack the U.S. govt.https://t.co/"
jenniferrenaud4|Moo57556470|-0.4943|0.2|0.714|0.086|"RT @Moo57556470: If Americans cannot trust its Congress, its FBI &amp; certainly its PEOTUS, how can we repair the damages absent A NEW ELECTIO"
cosmokramerss|MelindaThinker|0.2023|0.0|0.833|0.167|RT @MelindaThinker: Russian interference with the election could give courts legal authority to install Hillary https://t.co/By58AeeOe3
cosmokramerss|huffingtonpost|0.2023|0.0|0.833|0.167|RT @MelindaThinker: Russian interference with the election could give courts legal authority to install Hillary https://t.co/By58AeeOe3
ricknelms|summerbrennan|-0.4767|0.163|0.837|0.0|"RT @summerbrennan: As I've said before, I called McCain and Graham offices multiple times in tears right after the election and they are no"
BonnieSue05060|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
Tracy_Mack|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: @RandPaul just called for a bipartisan investigation into the issue of Russia messing with our election.Rand is a stand
eyetotelescope|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
bellablue1060|Green_Footballs|0.25|0.1|0.72|0.18|RT @Green_Footballs: One thing was confirmed beyond any doubt in this election: the Republican Party is just fine with white supremacism.
wmhsdemocrats|sethmoulton|0.6808|0.0|0.811|0.189|"RT @sethmoulton: Proud to see so many #MA6 constituents ready to work for change. There is so much to do, and this election was a call to a"
lucipujean|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
RobinWood|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
mcleans4|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
PageRemmers|Amy_Siskind|-0.4767|0.129|0.871|0.0|"RT @Amy_Siskind: When every poll, prognosticator and pundit is wrong on Election Night, and you say to yourself: how can this be?#russianh"
marilynmaupin|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
MarieMurcelle1|Pinkcloud15|0.2225|0.0|0.914|0.086|RT @Pinkcloud15: It's time 2 take our country back! Call the W H 202-456-1414 'n tell thm U want a new election done w/paper ballots! https
georgezab|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Yaznaa|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
JimW_JimW|breitbart|-0.296|0.128|0.872|0.0|Dem Sen McCaskill: Russian Involvement in Election a Form of Warfare - How breeds these fucking idiots https://t.co/TPf4AMxScT
AndyRichter|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
former_gop|amjoyshow|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
former_gop|t|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
facingdownfears|teenvogue|-0.1779|0.116|0.884|0.0|The BIG Way the Election Is Affecting People Who Have Anxiety #facingdownfears https://t.co/rJGAg1C9hE https://t.co/ok3zCQvTkJ
Pam24_CAbi|FaceTheNation|-0.0516|0.112|0.784|0.104|"RT @FaceTheNation: ""Russia tried to turn the election ... It means that Russia attacked the United States."" @TIME's Michael Duffy on CIA in"
TraceyRyniec|lazer_t|-0.4019|0.124|0.876|0.0|@lazer_t Investors in the railcar have been ignoring earnings for months. It wasn't just the Trump election. They're in denial.
PrettyBeaches|PattyMurray|0.3182|0.0|0.905|0.095|RT @PattyMurray: An investigation must begin as soon as possible on any evidence Russia actively worked to hijack our election &amp; elect Dona
pepperkatw|sallykohn|0.8495|0.0|0.646|0.354|"RT @sallykohn: If Russia had helped CLINTON win, can you imagine the GOP just quietly accepting it?!?!?!?https://t.co/57akQAyTrS"
pepperkatw|cnn|0.8495|0.0|0.646|0.354|"RT @sallykohn: If Russia had helped CLINTON win, can you imagine the GOP just quietly accepting it?!?!?!?https://t.co/57akQAyTrS"
george_gone|nathan2s1|-0.5473|0.227|0.773|0.0|RT @nathan2s1: MORE THAN HALF OF DETROIT'S VOTE-COUNTING MACHINES BROKE ON ELECTION DAYhttps://t.co/n8zQ33lQ4a
FLOURNOYFarrell|VampKiraLynn|0.3744|0.116|0.696|0.188|"@VampKiraLynn @retrosher @funder knowing again that the RUSSIAN government had rigged the election so he could win,"
Janie_St_K|_Makada_|-0.8074|0.307|0.693|0.0|RT @_Makada_: The same fake news media who said it was impossible to rig the election are now claiming Russia rigged the election with no p
itsjenlawrence|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
DebraMMason1|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
DebraMMason1|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
SoCalBIGmike|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
mtighe15|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
mtighe15|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
Ruthperricone|jamesplake721|-0.7555|0.244|0.756|0.0|RT @jamesplake721: CIA SAYS THE RUSSIANS GAVE THE ACTUAL VOTES TO @REALDONALDTRUMP #FAKENEWS AND ST UP LIES TO UNDERMINE THE ELECTION. DISG
DesignerDeb3|RealAlexJones|-0.7865|0.348|0.652|0.0|RT @RealAlexJones: #CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia - https://t.co/eXe3mPaIEG #infowars
DesignerDeb3|youtube|-0.7865|0.348|0.652|0.0|RT @RealAlexJones: #CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia - https://t.co/eXe3mPaIEG #infowars
1lisbongirl|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
BerkieBrenda|JasonLeopold|0.296|0.0|0.885|0.115|"RT @JasonLeopold: Key GOP senators join call for bipartisan Russia election probe, even as their leaders remain mumhttps://t.co/e1kISeZpap"
alexanderchee|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
DonnaMBaker3|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
travel611|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
travel611|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/FhGc6yE0ZI https://
RobMalara|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
magicalplatipus|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
magicalplatipus||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
cosmokramerss|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Just4Americans|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
redmcgraw1|tgreene319|0.0|0.0|1.0|0.0|RT @tgreene319: Let's review. CIA says Russian hackers interfered w election. Russia says they didn't. Trump doesn't believe CIA &amp; instead
Anyshka|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
NoveleraSalvaje|toddstarnes|0.8428|0.084|0.543|0.373|"RT @toddstarnes: Crowd:  Lock her up! Trump: That plays great before the election, now we dont care, right? Spoken like a true politic"
MarkingAround|DannyZuker|0.7184|0.0|0.76|0.24|"RT @DannyZuker: PATRIOT TEST:  If you're cool with Russia meddling with our election because your candidate won, you're not a patriot. Also"
trishforsythvos|cnn|0.5461|0.0|0.694|0.306|"I AGREE, bur how can we guard against cyber-hacking?! https://t.co/Nqo8v6YnSH"
bonniemac52|BryanDawsonUSA|-0.3612|0.135|0.865|0.0|RT @BryanDawsonUSA: GOP Congress:Hearings on #Benghazi witch hunt: 33Hearings on real Russian interference in US election: 0#russianha
inusanewscom|inusanews|0.5574|0.0|0.795|0.205|(Cbslocal) #Rep. #Moulton Tries To Foster Positive Response To Trump Election : It was.. https://t.co/rLXVXAXmBc https://t.co/71bxQcRUl4
BethAshworth5|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
rogiloc|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
marcylauren|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
marcylauren|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
goodtimenations|goodtimenation|-0.3182|0.15|0.85|0.0|Rajinikanths Said #Jayalalithaa Lost 1996 Tamil Nadu election because of me: South Indian https://t.co/xZIMOqJuBS
Kat4Obama|matthewamiller|-0.5106|0.202|0.798|0.0|RT @matthewamiller: Hard to miss the implication that Trump is going to put people in the IC to quash findings he disagrees with. https://t
Kat4Obama||-0.5106|0.202|0.798|0.0|RT @matthewamiller: Hard to miss the implication that Trump is going to put people in the IC to quash findings he disagrees with. https://t
Spartans4GOP|SenatorLankford|0.0|0.0|1.0|0.0|RT @SenatorLankford: TUNE IN: I'll be on Fox News tonight around 6:15pm ET to discuss Russian interference in the election. #russianhacking
AvieAvie47|claudiawrites|0.2187|0.109|0.743|0.147|RT @claudiawrites: Don't betray those who gave their lives fighting for their country. Investigate Russian ties to election. #CountryOverPa
marialenaj|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
deannawds|occupydemocrats|-0.1779|0.211|0.621|0.168|"POLITIFACT: Trump Is Lying, Russia DID Swing Election In His Favor - https://t.co/NskQ8X8Vac"
CriswellsOk|slone|0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
CriswellsOk||0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
blaha_b|abuhena0044|-0.1531|0.144|0.693|0.163|RT @abuhena0044: @HamiltonElector _Trump hijacked the election with Russian intervention committing treason to serve multiple interests at
CaroleBelew|mtracey|-0.25|0.095|0.905|0.0|"RT @mtracey: Dems' post-election lunacy closely resembles GOP birtherism, except in this case the paranoia is far more mainstream https://t"
CaroleBelew||-0.25|0.095|0.905|0.0|"RT @mtracey: Dems' post-election lunacy closely resembles GOP birtherism, except in this case the paranoia is far more mainstream https://t"
Heisse13|20committee|0.2023|0.0|0.924|0.076|RT @20committee: Trump's refusal to admit that Russia was behind election games is forcing his cabinet nominees to lie publicly in ways the
paul_carilli|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
paul_carilli|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
Yombe|2crazy4books2|0.0|0.0|1.0|0.0|RT @2crazy4books2: @Serpentine202 The CIA has proof. GOP conspired to suppress. https://t.co/UriwbWI930
Yombe|petitions|0.0|0.0|1.0|0.0|RT @2crazy4books2: @Serpentine202 The CIA has proof. GOP conspired to suppress. https://t.co/UriwbWI930
AliciaGs_BigMa|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
thecarlos3ff3ct|YouTube|0.296|0.104|0.714|0.182|"I liked a @YouTube video https://t.co/hRJsnlMQPV Morning Joe Host: Hillary Censored Us, Interfered In Election"
thecarlos3ff3ct|youtube|0.296|0.104|0.714|0.182|"I liked a @YouTube video https://t.co/hRJsnlMQPV Morning Joe Host: Hillary Censored Us, Interfered In Election"
Snap_Politics|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
Snap_Politics|t|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
DesignerDeb3|RealAlexJones|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
DesignerDeb3|infowars|-0.561|0.232|0.768|0.0|RT @RealAlexJones: MAXIMUM EMERGENCY! Rogue CIA Plans To Assassinate Trump Before Election - https://t.co/B0RXajXeLV
Lyn_Samuels|twitter|0.0|0.0|1.0|0.0|"Halt the election, EC and inauguration until we have a complete investigation of Russia, voting irregularities. https://t.co/5uGz4vJeGT"
ZangrawNOrlando|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
metamemette|metamemette|0.0|0.0|1.0|0.0|"RT @metamemette: @sethmoulton Let's see this in every Dem constituency in country, every month until the midterms. The election isn't over."
Ryan_Skalsky|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
taratemima|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
KarlaTKO|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
FlyingYogini|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
voilarie85210|voilarie85210|-0.25|0.136|0.777|0.087|RT @voilarie85210: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/Bashv9JORn via @P
voilarie85210|palmerreport|-0.25|0.136|0.777|0.087|RT @voilarie85210: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/Bashv9JORn via @P
TrumpismBook|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
gaylonparsons|Shoq|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
gaylonparsons|t|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
JoshuaCaseyGre2|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
simplyhoran|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
edgeoforever|ericgarland|-0.4404|0.116|0.884|0.0|"RT @ericgarland: But from about 2009 to the 2016 election, a madness is being brewed and slowly poured down the throats of increasingly hys"
Tracy_Mack|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
TheGOPJesus|feministabulous|0.0|0.0|1.0|0.0|RT @feministabulous: i can't believe russia would hack the election after trump specifically asked them to https://t.co/V1dTFKOZOa
TheGOPJesus|twitter|0.0|0.0|1.0|0.0|RT @feministabulous: i can't believe russia would hack the election after trump specifically asked them to https://t.co/V1dTFKOZOa
CEDADebate|cedadebate|0.7345|0.0|0.733|0.267|"The election results are in, thank you to everyone who ran and congrats to everyone who was elected!... https://t.co/nh5AFXLiZu"
e_revolutionist|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
e_revolutionist||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
ShadowClawDylan|aspen_eyes|0.5171|0.111|0.661|0.227|RT @aspen_eyes: GOD I'm so tired lmfaoForeign interference should invalidate an election. Period. But people seem all too happy to act li
bruleigh|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
bruleigh|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
DoorWay2Fandom|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
DoorWay2Fandom||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
MarieMurcelle1|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
shutupKatelynn|PolitiFact|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
shutupKatelynn|t|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
formarrowdbs|RepublicanChick|-0.1779|0.082|0.918|0.0|"RT @RepublicanChick: Liberals are accusing Russia of influencing the election. At the same time, liberals enabled citizens of other countri"
SandyTomich|summerbrennan|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
SandyTomich|t|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
Ravenchansan|ABCPolitics|0.0|0.0|1.0|0.0|RT @ABCPolitics: NEW: Bipartisan group of senators release joint statement calling for examination of reports of Russian interference in 20
ChrisGaryL|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
shrekandpearl|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
mmbaconomnom|JYSexton|-0.7003|0.264|0.652|0.084|RT @JYSexton: And for what? The election of a man who disgusts them and makes a mockery of their party. What a sad sack of shills these peo
linloy|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
linloy|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
jjsattorney|An0nKn0wledge|-0.6739|0.171|0.829|0.0|RT @An0nKn0wledge: THERE IS MORE EVIDENCE OF ALIENS EXISTING THEN THE RUSSIANS HACKING THE ELECTION.. BTW THE ELECTION FRAUD SO FAR ALL IN
realdadinstands|laurahollis61|-0.6486|0.238|0.762|0.0|"RT @laurahollis61: This whole ""Russians hacked the election"" story is the biggest load of crap since#Benghazi ""it-was-a-video."" Dems are d"
meltongoodwin|JohnWDean|0.0|0.0|1.0|0.0|RT @JohnWDean: The intel report on Russia's role in the 2016 election must be available for all electors before the electoral college meets
JanetETennessee|summerbrennan|-0.4767|0.163|0.837|0.0|"RT @summerbrennan: As I've said before, I called McCain and Graham offices multiple times in tears right after the election and they are no"
danielsofer|davewiner|-0.7579|0.279|0.636|0.085|"RT @davewiner: While we're outraged at Russian involvement in the election, the Repubs in Congress are killing Social Security, Medicare an"
paintedoctopus|RepFitzpatrick|0.296|0.0|0.864|0.136|@RepFitzpatrick Join the bipartisan effort 2 investigate #RussiaHacking If proven the election should b declared illegitimate #Putinspuppet
pmcnally202|KellyannePolls|0.3182|0.243|0.473|0.284|"@KellyannePolls there's a reason Duma broke into applause when he won election.  They know he weakens America, can be manipulated like child"
stksans|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
corygoings|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
TananariveDue|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
tericento|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
santiamtwit|twitter|-0.4767|0.193|0.807|0.0|Look who behind the Russian Fake News about Russian interference with election #maga https://t.co/bwZvRT6GTf
Th2shay|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Th2shay|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
rerrington1|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
MuseLotus|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
bakovic_steven|BryanDawsonUSA|-0.3612|0.135|0.865|0.0|RT @BryanDawsonUSA: GOP Congress:Hearings on #Benghazi witch hunt: 33Hearings on real Russian interference in US election: 0#russianha
wtflanksteak|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
wtflanksteak|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
today_global|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/wipAcVV1OV
laceylynn78|KeithOlbermann|-0.2023|0.139|0.75|0.111|"RT @KeithOlbermann: The Russians interfering in our election is, flatly, an act of war. From 9/28: is @realDonaldTrump loyal to the USA? ht"
sk8cello|DannyZuker|0.7184|0.0|0.76|0.24|"RT @DannyZuker: PATRIOT TEST:  If you're cool with Russia meddling with our election because your candidate won, you're not a patriot. Also"
simplyhoran|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
DavidJones2898|latimes|-0.0258|0.144|0.719|0.138|RT @latimes: Prominent senators say Russian election interference should alarm all Americans https://t.co/5QprDsvyoi https://t.co/SuFzJ25R0b
DavidJones2898|latimes|-0.0258|0.144|0.719|0.138|RT @latimes: Prominent senators say Russian election interference should alarm all Americans https://t.co/5QprDsvyoi https://t.co/SuFzJ25R0b
SuperPrivateEye|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
SoonerBeerSnob|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
Nomawrites|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
Purrpatrol|CarmineZozzora|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
Purrpatrol|t|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
pgcpro|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
pgcpro|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
SurfaceUnits|PrisonPlanet|-0.4939|0.276|0.724|0.0|@PrisonPlanet There is no evidence of any election hacking; let alone Russian hacking
maryaddie100|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
intenseCA|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Amy_Meeks|birbigs|-0.0387|0.05|0.95|0.0|RT @birbigs: There's evidence that Russia swayed the U.S. election &amp; we're supposed to NOT talk about it constantly? I'm sorry but that's u
1lisbongirl|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
rachelsYLG|freep|-0.4019|0.184|0.816|0.0|"Election day problems in MI ""one close election from a complete meltdown."" https://t.co/HxHAXP4Zg6 #AuditTheElection"
ladykayaker|DeanCathar|0.0|0.0|1.0|0.0|RT @DeanCathar: Send #CheetoLurch to jail BEFORE and the election becomes invalid#Theresistance#NotMyPresident@cspanwj https://t.co/hAX6
ladykayaker|t|0.0|0.0|1.0|0.0|RT @DeanCathar: Send #CheetoLurch to jail BEFORE and the election becomes invalid#Theresistance#NotMyPresident@cspanwj https://t.co/hAX6
dreece1480|MMFlint|0.8689|0.077|0.568|0.355|RT @MMFlint: The CIA has determined Russia hacked into our election to help elect Donald J. Trump. Now Trump names Putin best friend as OUR
davidhillgm|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
RanaeMayle|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
RanaeMayle|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
AaronMcCright|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
bsmart2b|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
bsmart2b|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
jumboglo|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
lorenz_louise|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
pattigandolfini|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
pattigandolfini|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
linloy|BryonWine|0.3182|0.066|0.806|0.128|"RT @BryonWine: McCain, Graham, Reed and Schumer questioning possible Russian influence in the election. Four Democrats. Yes, all DEMOCRATS."
fbrown7628|neeratanden|-0.636|0.257|0.743|0.0|@neeratanden @EricLiptonNYT @ScottShaneNYT @EricLichtblau everything is a ref to election! Who pays u to b depressing and loss of reality?
LynneAvVer|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
franksnstein|BruceBartlett|0.0|0.0|1.0|0.0|"RT @BruceBartlett: The question isn't why Russia interfered in our election, the question is why did in interfere on behalf of Trump &amp; the"
daletheamerica1|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Our favourite #FakeNews of the 2016 election https://t.co/Onm82JGBbn
daletheamerica1|twitter|0.0|0.0|1.0|0.0|RT @wikileaks: Our favourite #FakeNews of the 2016 election https://t.co/Onm82JGBbn
saintwalker98|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
BadCharacter77|hectormorenco|0.0|0.0|1.0|0.0|RT @hectormorenco: REAL NEWS: CIA &amp; MSM Make Up False Allegations of Russian Election Tampering Without Evidencehttps://t.co/jEyE0fR09S -
HeatherMoAndCo|ZaibatsuNews|0.2023|0.0|0.904|0.096|RT @ZaibatsuNews: WATCH: Chuck Todd hammers Reince Priebus over refusal to admit Russians might have influenced election https://t.co/ZuFWJ
HeatherMoAndCo|t|0.2023|0.0|0.904|0.096|RT @ZaibatsuNews: WATCH: Chuck Todd hammers Reince Priebus over refusal to admit Russians might have influenced election https://t.co/ZuFWJ
pugewok|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
pugewok|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
ggbootsrock|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
ggbootsrock|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
classygal21|TrumpsNewsDaily|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
classygal21|yahoo|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
JeffEKahn|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
JeffEKahn||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
DonnaVishio|JasonKander|-0.6597|0.213|0.787|0.0|"RT @JasonKander: If we ignore Russian espionage in our election, we embolden other foreign powers to launch similar attacks on every aspect"
sylvialyons981|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
Vuraelo_Reborn|kel12121|0.1531|0.178|0.581|0.24|RT @kel12121: I need to be like my dog he happy as hell the election didn't effect him. https://t.co/GOTVVgYgMY
Vuraelo_Reborn|twitter|0.1531|0.178|0.581|0.24|RT @kel12121: I need to be like my dog he happy as hell the election didn't effect him. https://t.co/GOTVVgYgMY
NIQUE_BELLA|joanneprada|-0.5719|0.381|0.619|0.0|RT @joanneprada: 2016 election: the ultimate scam
j3fk|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
j3fk|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
BlauesAugeBlond|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
otono60|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: BREAKING: Harry Reid says FBI Director James Comey deliberately withheld info on Russia's election meddling &amp; should re
MVkevinb|PrisonPlanet|-0.3453|0.139|0.861|0.0|RT @PrisonPlanet: Russia interfered in the election! (no evidence).LEFT FREAKS OUT.Saudi Arabia provably bankrolled Clinton's campaign.
laceylynn78|KeithOlbermann|0.0|0.0|1.0|0.0|"RT @KeithOlbermann: This was not an election, this was a Coup D'Etat abetted by traitors. From 11/1: The Trumpchurian Candidate https://t.c"
laceylynn78||0.0|0.0|1.0|0.0|"RT @KeithOlbermann: This was not an election, this was a Coup D'Etat abetted by traitors. From 11/1: The Trumpchurian Candidate https://t.c"
Veej_1|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
convoice|jahimes|0.0|0.0|1.0|0.0|@jahimes the people unhinged are those expecting the EC to reverse an election. Crybabies.
RickyLeeSongs|vicenews|-0.6808|0.259|0.741|0.0|"Here's a warning back in August. ""A foreign power could hack the US election, experts fear"" https://t.co/rUGbKUlETg via @vicenews"
RickyLeeSongs|news|-0.6808|0.259|0.741|0.0|"Here's a warning back in August. ""A foreign power could hack the US election, experts fear"" https://t.co/rUGbKUlETg via @vicenews"
monicasloves|politicususa|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
monicasloves|twitter|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
lgoldrick25|greenhousenyt|-0.0516|0.11|0.787|0.102|"RT @greenhousenyt: ""The fact that 59% of the vote-counting machines in Detroit all broke on Nov. 8 stands out as a stunning developmnt"" htt"
jdbashore|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
rhanser|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
rhanser|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
rphawg3150|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Mike_EH_52|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
mtighe15|davebernstein|-0.4019|0.114|0.886|0.0|RT @davebernstein: Former CIA agent Robert Baer said any other country would hold a new election they found out they were hacked. (6/10)htt
mrsperfectttt|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
alavecchia1|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
VPofClowns|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
hfsav001|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
SandiChilds|TwitterMoments|0.4588|0.063|0.75|0.188|RT @TwitterMoments: Top senators from both parties are banding together to demand an investigation into Russia's effect on the election. ht
DPMcCallum|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
dima7b_|twitter|-0.6249|0.203|0.797|0.0|"Mitch McConnell's role in this election is tantamount to treason. There is no way around this. What he did, was for https://t.co/dweCheTh8p"
huey_pat|LindaSuhler|-0.2168|0.144|0.75|0.106|RT @LindaSuhler: Remember Obama's hot mic msg to Putin about flexibility after the election?What are they scared of? #RussianHackinghttps
whatsmacksaid|thehighsign|-0.1027|0.065|0.935|0.0|RT @thehighsign: If only someone had tried to warn us about this Russian hacking business _before_the election. At a podium. During a debat
Trump4Pres0225|POTUSwas|-0.5106|0.163|0.837|0.0|.@POTUSwas given Morning briefs on CIA concerns with Russia involvement PRE ELECTION.  Where was the outrage THEN? https://t.co/nEpvwVX4rn
Trump4Pres0225|twitter|-0.5106|0.163|0.837|0.0|.@POTUSwas given Morning briefs on CIA concerns with Russia involvement PRE ELECTION.  Where was the outrage THEN? https://t.co/nEpvwVX4rn
alton_kalgae|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
thomasjoscelyn|jabeale|0.4019|0.0|0.881|0.119|"RT @jabeale: If Russia clandestinely interfered with a US election in order to favor a particular candidate, POTUS and the CIA should make"
Shawn22782896|PrisonPlanet|-0.3453|0.139|0.861|0.0|RT @PrisonPlanet: Russia interfered in the election! (no evidence).LEFT FREAKS OUT.Saudi Arabia provably bankrolled Clinton's campaign.
MARGARETFlana18|FiveRights|0.4215|0.094|0.697|0.209|"RT @FiveRights: Dear LiberalsThere was an election.You lost be bc you nominated a criminal.Rather than acting like 3rd world animals, tr"
deanrcarey|wikileaks|-0.1027|0.122|0.778|0.1|RT @wikileaks: Police admit sex complaint against Assange was fabricated in elaborate plot https://t.co/OPCFRveUqM More: https://t.co/Mb6gX
deanrcarey|mcclatchydc|-0.1027|0.122|0.778|0.1|RT @wikileaks: Police admit sex complaint against Assange was fabricated in elaborate plot https://t.co/OPCFRveUqM More: https://t.co/Mb6gX
riledirish|KeepAmerGr8|-0.5719|0.222|0.778|0.0|RT @KeepAmerGr8: Bipartisan anger grows over Russian interference into U.S. election https://t.co/9MgHpkwma0 via @HuffPostPol
riledirish|huffingtonpost|-0.5719|0.222|0.778|0.0|RT @KeepAmerGr8: Bipartisan anger grows over Russian interference into U.S. election https://t.co/9MgHpkwma0 via @HuffPostPol
KenBerry611|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
KenBerry611|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
ThatLaddChick|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
HindmanDebra|BreitbartNews|-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
HindmanDebra||-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
BevPerryMusic|EricBoehlert|0.0|0.0|1.0|0.0|"RT @EricBoehlert: this is why, to date, we have to rely on anonymous sources for information re: Russia and election https://t.co/OSbrbw66M5"
BevPerryMusic|twitter|0.0|0.0|1.0|0.0|"RT @EricBoehlert: this is why, to date, we have to rely on anonymous sources for information re: Russia and election https://t.co/OSbrbw66M5"
JoeMacPhail|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
lifeandstuff247|FitzyGFY|-0.7574|0.319|0.681|0.0|RT @FitzyGFY: I'm w/@mtdisme - Russia absolutely hacked into Steelers PSI last week to distract from US election accusations #DeflateGate2
BrownGig|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
AndreLinoge68|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
tonecky|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
StoneColdChik|icowrich|-0.6239|0.267|0.733|0.0|"@icowrich @nytimes right, before hilary lost the election she thought she had rigged to the hilt!"
mkisswag|Holbornlolz|-0.6705|0.231|0.684|0.085|RT @Holbornlolz: People who killed 100's of 1000's to ensure regime change all over the M. East are upset that Russia may have interfered i
Shoepirate|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
pathogen43|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
ojhines2k|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
ojhines2k|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
NYtitanic1999|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
NYtitanic1999|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
veve4heart|TechCrunch|0.0|0.0|1.0|0.0|RT @TechCrunch: Obama orders review of Russian election hacking https://t.co/AF9SI1AMtU
veve4heart|techcrunch|0.0|0.0|1.0|0.0|RT @TechCrunch: Obama orders review of Russian election hacking https://t.co/AF9SI1AMtU
alavecchia1|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
KTynot|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
tlhenson823|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
USNCS|ShortCanuck|-0.5719|0.188|0.812|0.0|@ShortCanuck @summerofsoaps @mermaidaysh @yasmin86 @ghoulette27 I don't think I had chatted with her since the election. Man I hate that.
tadpoledrain|BrendanNyhan|-0.4659|0.169|0.787|0.043|"RT @BrendanNyhan: Seeing people dismiss as silly conspiracy talk, but far more serious. Potential Dep SOS suggesting Obama used IC in a dom"
edenfan|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Other than @LindseyGrahamSC is there a single principled Republican in Washigton? Russia directly intervened in our electio
JanFrye|americanthinker|0.4215|0.0|0.741|0.259|Blog: Obama's CIA: Russians favored Trump in election https://t.co/in6U9kQdYm
Ghifarix|ggreenwald|0.4471|0.075|0.774|0.15|RT @ggreenwald: The combination of Corbyn &amp; Brexit sent the UK political/media class into sustained madness but it's nothing compared to po
SovietGuacamole|twitter|-0.4767|0.134|0.866|0.0|Black women have always been historically deprived of their rights. Why did it take this election to realize how mu https://t.co/KTqgDP5D3r
indee2|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
thednaofmath|12voltman60|0.2944|0.0|0.901|0.099|"RT @12voltman60: @FoxNews @WTPatty @JudgeJeanine Remember his ""hot mic"" moment in '12 with Russia saying he'd be more flexible after the e"
mateosfo|anirvan|0.6486|0.0|0.806|0.194|"RT @anirvan: Huge props to 50+ stores across #Berkeley, CA that put up ""Everyone is Welcome Here"" posters, in the wake of 14 post-election"
Nomawrites|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
iru_guy|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
pgrandee10|HuffingtonPost|0.0|0.0|1.0|0.0|RT @HuffingtonPost: Trump pays his own businesses $3 million in days surrounding election https://t.co/ng40HjL3ur https://t.co/PaFNg7vAdF
pgrandee10|m|0.0|0.0|1.0|0.0|RT @HuffingtonPost: Trump pays his own businesses $3 million in days surrounding election https://t.co/ng40HjL3ur https://t.co/PaFNg7vAdF
mslizag|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
metamemette|sethmoulton|0.0|0.0|1.0|0.0|"@sethmoulton Let's see this in every Dem constituency in country, every month until the midterms. The election isn't over. #Win2018 #mapoli"
AlexHSTL|tomtomorrow|-0.7841|0.247|0.703|0.05|RT @tomtomorrow: Thought of what Trump's election means for this country has left me feeling the sort of grief I have felt after death of s
Model41081|scottwongDC|-0.34|0.112|0.888|0.0|"RT @scottwongDC: In rare bipartisan statement, McCAIN, GRAHAM, SCHUMER &amp; REED say reports of Russian interference in election ""should alarm"
redmor11|Peter_Wehner|0.743|0.0|0.741|0.259|"RT @Peter_Wehner: Rs shrugging off Russian intervention in our election is a perfect illustration of what @JonHaidt refers to as ""motivate"
hamel1776|youtube|-0.1531|0.127|0.873|0.0|"Morning Joe Host: Hillary Censored Us, Interfered In Election https://t.co/B8pqAV5NFd #YouTube #TheAlexJonesChannel"
Kwayylo|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
GeNes1S21|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
dajosc11|timcarvell|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
dajosc11|freep|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
smartvalueblog|slone|0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
smartvalueblog||0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
RandyCFord|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
bkg713|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
sarat_varanasi|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
abhasharma61|GitRDoneLarry|0.7084|0.124|0.612|0.264|RT @GitRDoneLarry: I know I said I'm blocking all Whiney election tweet but some are so dad gum entertaining! Ok starting again... now.
aadisharma1900|TimesNow|-0.0366|0.176|0.659|0.165|@TimesNow Don't do that if u dont wanna lose the election shamelessly
sekairider|chucktodd|-0.3382|0.094|0.906|0.0|"If only the MSM &amp; @chucktodd knew about @HillaryClinton's email server during the election. I bet they'd get to the bottom of it! But, alas."
Fnwy|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
dougnot2|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
bikerbd|PolitixGal|-0.8519|0.364|0.636|0.0|RT @PolitixGal: DEMS &amp; Clintons are desperate to blame someone other than themselves for their election loss. Hillary was a liar who didn't
tsujigo|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
realmojesse5372|GartrellLinda|0.0|0.0|1.0|0.0|RT @GartrellLinda: Netanyahu pollsterObama role in election larger than reported https://t.co/ZiixnPXfbS HYPOCRITES interfered in Israeli e
realmojesse5372|thehill|0.0|0.0|1.0|0.0|RT @GartrellLinda: Netanyahu pollsterObama role in election larger than reported https://t.co/ZiixnPXfbS HYPOCRITES interfered in Israeli e
4TruthAndReason|poodbit499|-0.516|0.21|0.696|0.094|"RT @poodbit499: Yes OBAMA hates BiBi so much he interfered w/Israels election &amp; tried to oust him,yet he's trying 2 BLAME Russia 4 HRC bein"
LindaFrum|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
LindaFrum||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
JebCuck|BreitbartNews|-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
JebCuck||-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
KenicVerlene|WithCongress|-0.5267|0.167|0.833|0.0|"@WithCongress Rahul Stupid Donkey parliament is not your Mommy's property, next Election Public going to kick your https://t.co/udsH5FNRUA"
KenicVerlene|twitter|-0.5267|0.167|0.833|0.0|"@WithCongress Rahul Stupid Donkey parliament is not your Mommy's property, next Election Public going to kick your https://t.co/udsH5FNRUA"
tootropic|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
tootropic|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
AGMcThugabobs|An0nKn0wledge|-0.6739|0.171|0.829|0.0|RT @An0nKn0wledge: THERE IS MORE EVIDENCE OF ALIENS EXISTING THEN THE RUSSIANS HACKING THE ELECTION.. BTW THE ELECTION FRAUD SO FAR ALL IN
2lisa4|quinncy|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
2lisa4|palmerreport|-0.3612|0.122|0.878|0.0|"RT @quinncy: Rigged election: months ago, Steve Bannon ""knew"" precisely which states Donald Trump would flip https://t.co/F5KNTgdUj6 via @P"
WomanVote|laureldavilacpa|0.0|0.0|1.0|0.0|RT @laureldavilacpa: #ImStillNotOver Before the election the Senate was briefed by the CIA of #RussianHackers electioneering for Trump - an
Tracy_Mack|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
kmclc2016brutus|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
DKWilson56|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
DKWilson56|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
rphawg3150|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
buckycapped|DrGMLaTulippe|0.5927|0.0|0.851|0.149|"RT @DrGMLaTulippe: It'll take you ten minutes to read this thread, but it's imperative that you do.First thing that's made me feel better"
RalphHornsby|youtube|0.0|0.0|1.0|0.0|CIA Splinter Group Calls For Overthrow Of Trump Election - YouTube https://t.co/On5QWnznSl
jsim63|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
jsim63||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
ThomasBialek2|chuckwoolery|0.0|0.0|1.0|0.0|RT @chuckwoolery: Libs say #Trump stole the election but Dems actually handed it to him. @MarkYoungTruth explains on #BluntForceTruth https
M_CollinsDesign|HouseofCards|-0.2183|0.144|0.755|0.101|America was so impatient for new seasons of @HouseofCards and @VeepHBO that we created the 2016 election.
CuriousCat1950|twitter|0.8779|0.0|0.598|0.402|Election shows clearly many of t 'flaws' in US system in glorious Technicolor. Looking pretty Mickey Mouse. Remedie https://t.co/wpOakbh4xK
Cici0804|RisaWechsler|0.3182|0.0|0.905|0.095|"RT @RisaWechsler: If @leahmcelrath 's thread made you curious abt Dugin, watch what he had to say about election and its consequences. http"
bossclockwork|mrpcunningham|0.0|0.0|1.0|0.0|"RT @mrpcunningham: In modern Russia, election interferes with you!"
macvolley1|MissLizzyNJ|-0.952|0.53|0.47|0.0|"RT @MissLizzyNJ: #ImStillNotOver the fact that I lost the election because I'm a lying criminal and America hates me, so I'll blame fake ne"
jjmac818|ACNewman|0.34|0.124|0.659|0.217|"RT @ACNewman: Look, more shadiness in the election. If true, Michigan was stolen. If that's true, why not others ? https://t.co/OSorsOpmO0"
jjmac818|palmerreport|0.34|0.124|0.659|0.217|"RT @ACNewman: Look, more shadiness in the election. If true, Michigan was stolen. If that's true, why not others ? https://t.co/OSorsOpmO0"
DViper22|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
DViper22|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
EnigmaNetxx|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
EnigmaNetxx|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
amandelman|bamendelsohn|0.0|0.0|1.0|0.0|"@bamendelsohn 2 weeks ago, UW-Madison hosted a public panel re: the election, conducted as if not one of 200 ppl present was conservative"
Patta47cake|jahimes|0.6375|0.0|0.754|0.246|RT @jahimes: @GoodJobGuru @PoliticalLine Yes. The election is over. But the electoral college has not met. So no President has been legally
EzabQuader|LOLGOP|0.25|0.058|0.846|0.096|RT @LOLGOP: This election is like if A Christmas Carol ended with Scrooge getting a giant tax break paid for by cutting Tiny Tim off Medica
_mommapie|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
LilRedheaad|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
AdamPacton|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
mtighe15|TomthunkitsMind|0.0|0.0|1.0|0.0|RT @TomthunkitsMind: Russia Says It Was In Touch With Trump Campaign During The Election. https://t.co/ik0yyqk7fF https://t.co/g7PF8uOlfg
mtighe15|huffingtonpost|0.0|0.0|1.0|0.0|RT @TomthunkitsMind: Russia Says It Was In Touch With Trump Campaign During The Election. https://t.co/ik0yyqk7fF https://t.co/g7PF8uOlfg
shaquita025|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
my_opinion_man|ABCPolitics|0.0|0.0|1.0|0.0|RT @ABCPolitics: NEW: Bipartisan group of senators release joint statement calling for examination of reports of Russian interference in 20
mmaureen7|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Mike_EH_52|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
blueinthesouth|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
blueinthesouth|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
Diamondrosegrfx|MadJewessWoman|0.0|0.0|1.0|0.0|"RT @MadJewessWoman: .@realDonaldTrumpINVESTIGATE @SenJohnMcCain 4 overthrowing #Ukraine govt, influencing election in #KIEV, 2013-14http"
bigbabe2022|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: BREAKING: Harry Reid says FBI Director James Comey deliberately withheld info on Russia's election meddling &amp; should re
penny63434309|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
penny63434309|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
AlgoENews|nypost|0.5859|0.0|0.759|0.241|How political rags reacted to Donald Trumps election win https://t.co/ATzE2bD6zz #enews #Trending https://t.co/FdE8sn0Aea
DeanCathar|cspanwj|0.0|0.0|1.0|0.0|Send #CheetoLurch to jail BEFORE and the election becomes invalid#Theresistance#NotMyPresident@cspanwj https://t.co/hAX6bMXMLi
DeanCathar|twitter|0.0|0.0|1.0|0.0|Send #CheetoLurch to jail BEFORE and the election becomes invalid#Theresistance#NotMyPresident@cspanwj https://t.co/hAX6bMXMLi
FashionHitList|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
Serabbi|SenatorTomUdall|0.5267|0.067|0.714|0.219|RT @SenatorTomUdall: I will join lawmakers in both parties &amp; demand investigation of Russia's effort to influence presidential election. ht
internet_dad69|JhonRules|-0.4019|0.124|0.876|0.0|"RT @JhonRules: date: can you believe russia hacked the u.s. to change the electionme, leaning in: i would never hack you"
Marie_Al_Marie|yahoo|0.0|0.0|1.0|0.0|"Watch what they do, don't listen to what sociopathic people say. https://t.co/k7aJj23W31"
KerryCounahan|ezlusztig|-0.0688|0.059|0.891|0.049|RT @ezlusztig: THE FBI STOLE THIS ELECTION. Don't forget it. And don't wake up tomorrow and decide you have no choice but to live with it.
SnowdenMark1|openquotes|0.0|0.0|1.0|0.0|"During the 2000 election, the current administration told our milit... #IkeSkelton #quotations https://t.co/iyHBFmGrLr"
TreyArline|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
VollmerAntes|emrutherford90|-0.5423|0.176|0.824|0.0|"RT @emrutherford90: Member when Russia forced H to set up a private server in home, rig the dem election, use BleachBit to erase. Then made"
asiannicensweet|NoceraNYT|0.0|0.0|1.0|0.0|RT @NoceraNYT: Is this for real?  https://t.co/AHODO2pTpa
asiannicensweet|palmerreport|0.0|0.0|1.0|0.0|RT @NoceraNYT: Is this for real?  https://t.co/AHODO2pTpa
ubervaper|tgreene319|0.0|0.0|1.0|0.0|RT @tgreene319: Let's review. CIA says Russian hackers interfered w election. Russia says they didn't. Trump doesn't believe CIA &amp; instead
peacelovedixie|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
julianwilson38|BardockObama|-0.8208|0.322|0.591|0.087|"RT @BardockObama: Liberals are so stupid y'all ask for a recount then fail, then think Russia rigged the election lol it was obviously J Co"
dleeprice|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
dleeprice|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
knowlton_paula|ezlusztig|0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
knowlton_paula||0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
Landwehr_Erik|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
adamlparker|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
adamlparker|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
smell3roses|JasonLeopold|0.296|0.0|0.885|0.115|"RT @JasonLeopold: Key GOP senators join call for bipartisan Russia election probe, even as their leaders remain mumhttps://t.co/e1kISeZpap"
KarrenKuk|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
chavezglen1755|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/mEIzELKuVz https://t."
chavezglen1755||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/mEIzELKuVz https://t."
DestructiveChem|DavidAFrench|-0.3612|0.122|0.878|0.0|RT @DavidAFrench: What's the argument against a bipartisan investigation of Russian efforts to disrupt and/or influence the election? Is th
trupatriot4|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
trupatriot4|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
ekangas81|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
Sharonsayswhat|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
IAmChey_D|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
IAmChey_D|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
sssssssssaamm|vicenews|-0.3612|0.116|0.884|0.0|"RT @vicenews: I think its ridiculous"" Trump continues to shrug off a CIA report that Russia meddled in the 2016 election https://t.co/p6m"
sssssssssaamm|t|-0.3612|0.116|0.884|0.0|"RT @vicenews: I think its ridiculous"" Trump continues to shrug off a CIA report that Russia meddled in the 2016 election https://t.co/p6m"
plbrocks|Vassa42|-0.4019|0.109|0.891|0.0|RT @Vassa42: It is widely expected that Daniel Andrews &amp; his disaterois Labor Govt will lose the 2018 Vic State Election. #springst https:/
plbrocks||-0.4019|0.109|0.891|0.0|RT @Vassa42: It is widely expected that Daniel Andrews &amp; his disaterois Labor Govt will lose the 2018 Vic State Election. #springst https:/
RobinBall1961|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
nakhon224|tass|0.5267|0.0|0.673|0.327|"""Legislature speaker winning presidential election in Moldovas"" https://t.co/YaCWC8fkgJ"
Stopcnnlies|hautedamn|-0.34|0.113|0.833|0.054|RT @hautedamn: The people who want you to believe Russia hacked the election are the same people telling you #pizzagate isn't real.
WVIndependent|PolitiFact|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
WVIndependent|t|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
edenfan|GeorgeTakei|0.0|0.0|1.0|0.0|"RT @GeorgeTakei: The CIA assessment concludes that Russians interfered with our election. With the margin so close, the result is illegitim"
575haiku|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
IamHer847|North_Socialist|0.0|0.0|1.0|0.0|@North_Socialist And he knew about the infiltration and still released the letter one week before the election. Hmmm!
MarkopoloXYZ|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
MarkopoloXYZ|change|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
Donny160170|veggie64_leslie|-0.3016|0.145|0.759|0.096|"RT @veggie64_leslie: Homeland Security IP address linked to attempted hack into GA voting systemIs this ""fake news"" HRC was afraid of?htt"
getrealvonciel|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
getrealvonciel|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
Pyt2008Yvonne|emigre80|-0.3802|0.217|0.662|0.121|"RT @emigre80: Both Trump and Sanders were delighted to cry ""rigged election!"" when they ran against Clinton.Now that there's evidence? *C"
juneday864|casatino|-0.1027|0.097|0.903|0.0|RT @casatino: FBI: sends vague letter; actually nothingMSM: *quivers*CIA: confirms Russia interfered w/electionMSM: \_()_/https://
mr_dsantos|TeaPainUSA|-0.4215|0.141|0.859|0.0|"RT @TeaPainUSA: This is the first election in American history that the incoming President is the ""lame duck."""
FLOURNOYFarrell|VampKiraLynn|-0.3612|0.106|0.894|0.0|@VampKiraLynn @retrosher @funder several systems and later he tried to cover telling on himself by saying that the election system is rigged
INVUQT|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: What if the election hadn't been hacked?What if Hillary hadn't stole the nomination?What if Obama hadn't given rise to
adellelalane|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/oinoIzHBra
butzmom|DavidCornDC|-0.5095|0.272|0.623|0.105|"@DavidCornDC ""Outrage"" is a bit misleading. More preventing future cyber attacks of the parties than Russian attempt to sway 2016 election."
MaximusAthos|HuffPostPol|-0.5719|0.252|0.748|0.0|Bipartisan anger grows over Russian interference into U.S. election https://t.co/s60Sz4dFrH # via @HuffPostPol
MaximusAthos|huffingtonpost|-0.5719|0.252|0.748|0.0|Bipartisan anger grows over Russian interference into U.S. election https://t.co/s60Sz4dFrH # via @HuffPostPol
taurocephala|NPR|0.3612|0.0|0.848|0.152|Via @NPR: Reporter's Notebook: What It Was Like As A Muslim To Cover The Election https://t.co/Jx15CwT5Lp
taurocephala|npr|0.3612|0.0|0.848|0.152|Via @NPR: Reporter's Notebook: What It Was Like As A Muslim To Cover The Election https://t.co/Jx15CwT5Lp
ClaytonMuirhead|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Our favourite #FakeNews of the 2016 election https://t.co/Onm82JGBbn
ClaytonMuirhead|twitter|0.0|0.0|1.0|0.0|RT @wikileaks: Our favourite #FakeNews of the 2016 election https://t.co/Onm82JGBbn
ShanksTheAuthor|HartoshSinghBal|0.0772|0.235|0.504|0.261|@HartoshSinghBal The election rhetoric insults our intelligence so.
ladykayaker|MrBudSmith|0.2023|0.0|0.904|0.096|RT @MrBudSmith: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/8xo
ladykayaker|t|0.2023|0.0|0.904|0.096|RT @MrBudSmith: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/8xo
SwaggyP_803|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
SwaggyP_803|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
lizfdonohue|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
mainemama48|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
Tuffelhund2003|Meow1113|0.0|0.0|1.0|0.0|@Meow1113 4.8M petition signers aren't changing an election that 120M voted in.
vanduynje|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
sacpros|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/bJR3VATU5P
lynnguppy|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
DavenportIowaa|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/AZF8IyF2Oj #Davenport #Iowa
EbiGahama|2dJazz|0.7845|0.0|0.685|0.315|RT @2dJazz: Arc System Works Awards 2016 election results:GG: @koichinko &amp; @gou4th_fab BB: @soujif91 &amp; @MINAMI_IZANAMI Congratulations 
3rdrockhome|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/hehKt08KAT #TopStories
PaedoAbuseLiars|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News: Washington Post https://t.co/O4VvO0uNgO #TopStories #paedobritain
ploop52|emmartin173|0.6369|0.0|0.776|0.224|RT @emmartin173: @charles_gaba Qs: has MSM learned anything about Republicans since election? Do they know they normalized R Party like the
etalbert|PeterFosterALP|-0.4588|0.15|0.85|0.0|RT @PeterFosterALP: What a fizza.No wonder Australians are fed up with all the deceit of Malcolm Turnbulls fraudband https://t.co/ZEVqV
etalbert|t|-0.4588|0.15|0.85|0.0|RT @PeterFosterALP: What a fizza.No wonder Australians are fed up with all the deceit of Malcolm Turnbulls fraudband https://t.co/ZEVqV
kfpeters|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
StevenNantz|PattyMurray|0.6124|0.0|0.737|0.263|"@PattyMurray Yes. Senator, please insist on a bipartisan investigation of Russian intervention in the 2016 presidential election"
matt_spiro|ParkerMolloy|-0.5067|0.17|0.83|0.0|"RT @ParkerMolloy: ""patrioteagle.flag says there's a child sex pizza dungeon!""""On it!""""The CIA says Russia messed w/ the election!""Some s"
bonita_jay1|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
bonita_jay1|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Shepherdof9|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
EllenMorris1222|JoyAnnReid|0.0|0.0|1.0|0.0|"RT @JoyAnnReid: And by the way if @SenatorReid is right, and the head of the FBI stood by and let Russia meddle in our election (then did s"
silver_selkie|leahmcelrath|0.5584|0.0|0.796|0.204|RT @leahmcelrath: Watergate seems like such an minor almost innocent bit of subterfuge compared to what's happened in this election.
cbba21|Sifill_LDF|-0.5423|0.137|0.863|0.0|RT @Sifill_LDF: Everyone outraged by this foreign interference in our election should be on the phone 1st thing Mon to their Reps.  https:/
cbba21||-0.5423|0.137|0.863|0.0|RT @Sifill_LDF: Everyone outraged by this foreign interference in our election should be on the phone 1st thing Mon to their Reps.  https:/
BevPerryMusic|ProudlyLiberal2|-0.5994|0.17|0.83|0.0|"RT @ProudlyLiberal2: KeithOlbermann: The Russians interfering in our election is, flatly, an act of war. From 9/28: is realDonaldTrump  ht"
blueskymountain|MariefromPA|0.0|0.0|1.0|0.0|@MariefromPA everything in this election has been unprecedented &amp; since rules don't seem to apply anymore... who knows (??)
naenae_away|jenanne34|0.8176|0.0|0.653|0.347|"@jenanne34 ""Liberals"" really think the election of a huge diverse country like America should be won by only appeal https://t.co/TxcC0Qkag1"
naenae_away|twitter|0.8176|0.0|0.653|0.347|"@jenanne34 ""Liberals"" really think the election of a huge diverse country like America should be won by only appeal https://t.co/TxcC0Qkag1"
fatousaidykhan|Smith_JeffreyT|0.1531|0.122|0.732|0.146|RT @Smith_JeffreyT: RE: Jammeh taking election defeat to #Gambia's Supreme Court: hearing must happen w/in 10 days after election. Monday =
StarKat99|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
lawwtey|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
genericlogin|PolitiFact|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
genericlogin|t|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
mowapello604|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
guyinblackhat|medium|-0.1531|0.12|0.787|0.093|"""Russia manipulated our election and ... appear poised to install their puppet into the presidency of our nation."" https://t.co/1Cc00kfISb"
DeborahKayGilb2|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
DeborahKayGilb2|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
sarahtimmerman|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
walkileaks|walkileaks|0.0|0.0|1.0|0.0|Eric Shawn reports: The alleged Russian electionhacking https://t.co/3itAsmnpiX
DeniseJeffress|Franklin_Graham|-0.3182|0.113|0.887|0.0|RT @Franklin_Graham: The media were shocked by the real difference made by evangelical voters in the last election. https://t.co/6lUOVf96zA
DeniseJeffress|m|-0.3182|0.113|0.887|0.0|RT @Franklin_Graham: The media were shocked by the real difference made by evangelical voters in the last election. https://t.co/6lUOVf96zA
RandyCFord|fitness_linda|0.4215|0.0|0.797|0.203|@fitness_linda @thehuntinghouse @mtraceyLike your actions are to destabilize faith in the election?
d0g0fd0ggerland|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
d0g0fd0ggerland|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
MissKanuck|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
HighOnFloyd|voxdotcom|0.0|0.0|1.0|0.0|"Russia's role in this year's presidential election, explained by a media historian https://t.co/HkcVYrKII0 via @voxdotcom"
HighOnFloyd|vox|0.0|0.0|1.0|0.0|"Russia's role in this year's presidential election, explained by a media historian https://t.co/HkcVYrKII0 via @voxdotcom"
lalawatsup|VanJones68|0.6988|0.0|0.757|0.243|@VanJones68 Just saw your post election appearance on @TheDailyShow.  Thank you for upcoming special! don't give them all to trump!
BigSwingTheory|ericgarland|-0.4404|0.116|0.884|0.0|"RT @ericgarland: But from about 2009 to the 2016 election, a madness is being brewed and slowly poured down the throats of increasingly hys"
Coreybez1|FoxNews|-0.7783|0.466|0.46|0.075|"RT @FoxNews: Latest excuse - @HillaryClinton blames election loss on ""fake news."" https://t.co/UgjfIZUALc"
Coreybez1|twitter|-0.7783|0.466|0.46|0.075|"RT @FoxNews: Latest excuse - @HillaryClinton blames election loss on ""fake news."" https://t.co/UgjfIZUALc"
BJeanMohr1|amjoyshow|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
BJeanMohr1|t|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
Based_Gibson|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
niknamH|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
ElaineFox|ByronYork|0.0|0.0|1.0|0.0|RT @ByronYork: Vote totals in Mike Pence's DC neighborhood. 309 people in precinct voted Trump/Pence. Staying mostly quiet. https://t.co/3c
ElaineFox|t|0.0|0.0|1.0|0.0|RT @ByronYork: Vote totals in Mike Pence's DC neighborhood. 309 people in precinct voted Trump/Pence. Staying mostly quiet. https://t.co/3c
oxbeyedoc|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
oxbeyedoc|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
Woolndoghairs|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
xfigmentx|summerbrennan|-0.4767|0.163|0.837|0.0|"RT @summerbrennan: As I've said before, I called McCain and Graham offices multiple times in tears right after the election and they are no"
Ellesun|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
momof3moochers|JudgeJeanine|0.0|0.0|1.0|0.0|"RT @JudgeJeanine: ""The election is over - you're either with us or against us. That is...with the U.S. or against the U.S.""-@JudgeJeanine #"
LindaLeeJones11|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
Zanzan280|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/4TnN8g6MGt https://t."
Zanzan280||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/4TnN8g6MGt https://t."
WonderWinged|RBReich|0.3612|0.0|0.848|0.152|"@RBReich I think we should put the election and move on , it's like running in circle"
ChrisParry|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
AJeanRuggiero|ElectoralCollge|-0.4184|0.202|0.798|0.0|. @ElectoralCollge This in addition 2 colluding w/Russia to tamper election.TREASON! TREASON!@GOP @TheJusticeDept https://t.co/T6bVdDQt4Q
AJeanRuggiero|twitter|-0.4184|0.202|0.798|0.0|. @ElectoralCollge This in addition 2 colluding w/Russia to tamper election.TREASON! TREASON!@GOP @TheJusticeDept https://t.co/T6bVdDQt4Q
CYNJONES|DrBelasen|0.0|0.0|1.0|0.0|"RT @DrBelasen: @MissVociferous @JohnWDean Trump is compromised. Regardless of the status of the recount, the results of the election are fl"
h0tbreakingnews|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/1sdoYa4jvj #BreakingNews
guna15|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
guna15|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
PeteKaliner|DavidAFrench|-0.3612|0.122|0.878|0.0|RT @DavidAFrench: What's the argument against a bipartisan investigation of Russian efforts to disrupt and/or influence the election? Is th
nick_at_dev|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
magicalplatipus|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
withlovenao|EJjuninho|0.0|0.0|1.0|0.0|RT @EJjuninho: 10. Bernie Sanders would've washed Trump in the election.
VetApologist|SarahPalinUSA|-0.0422|0.118|0.77|0.112|RT @SarahPalinUSA: Russia's getting out of hand? So says the defeated. Not to worry... remember I can keep an eye on them from here. https:
LyndaPole|AnaCosentino2|-0.0772|0.199|0.664|0.137|RT @AnaCosentino2: @dissentingj @LyndaPole @CNBC @NBCNews No patience 4 Millennials..your protest vote handed election 2 Bozo.I hope you st
tleydn|chucktodd|0.7506|0.0|0.748|0.252|@chucktodd awesome job today grilling @Reince on whether he believes CIA assertion of Russian interference of US election. Please grill more
miltoncosta|PokitDok|0.0|0.0|1.0|0.0|RT @PokitDok: The election results are in and it could be a big change for the #ACA and future of healthcare. Learn why: https://t.co/44VBg
miltoncosta|t|0.0|0.0|1.0|0.0|RT @PokitDok: The election results are in and it could be a big change for the #ACA and future of healthcare. Learn why: https://t.co/44VBg
spzkaz|MissLizzyNJ|-0.952|0.53|0.47|0.0|"RT @MissLizzyNJ: #ImStillNotOver the fact that I lost the election because I'm a lying criminal and America hates me, so I'll blame fake ne"
emily_lombardi|feministabulous|0.0|0.0|1.0|0.0|RT @feministabulous: i can't believe russia would hack the election after trump specifically asked them to https://t.co/V1dTFKOZOa
emily_lombardi|twitter|0.0|0.0|1.0|0.0|RT @feministabulous: i can't believe russia would hack the election after trump specifically asked them to https://t.co/V1dTFKOZOa
ciardha|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
ciardha||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
WintersNFL|twitter|-0.2732|0.174|0.826|0.0|I'm still blocked by the zombie even after the election. https://t.co/XCKV4PxJRp
RIMURO|amjoyshow|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
RIMURO|t|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
speedyeproducts|chicagotribune|0.0|0.0|1.0|0.0|2) https://t.co/HDoiwJ0iwA
kmqkatie|ASquareOfSkye|0.0|0.0|1.0|0.0|RT @ASquareOfSkye: Russian-backed Paul Manafort told Donald Trump to target Michigan just before Election Day https://t.co/NWYB70Un2C via @
kmqkatie|palmerreport|0.0|0.0|1.0|0.0|RT @ASquareOfSkye: Russian-backed Paul Manafort told Donald Trump to target Michigan just before Election Day https://t.co/NWYB70Un2C via @
donaldwatkins01|ABC|-0.5826|0.166|0.834|0.0|@ABC @MLevineReports There is where they will find the method in the election result deception ! Keep looking! It is there!
bad_indian_girl|JasonKander|-0.6597|0.213|0.787|0.0|"RT @JasonKander: If we ignore Russian espionage in our election, we embolden other foreign powers to launch similar attacks on every aspect"
BoxANT|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
danmonaghan|summerbrennan|-0.4767|0.163|0.837|0.0|"RT @summerbrennan: As I've said before, I called McCain and Graham offices multiple times in tears right after the election and they are no"
N4LRB4me|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
N4LRB4me|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
quarklesparkle|MrBudSmith|0.2023|0.0|0.904|0.096|RT @MrBudSmith: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/8xo
quarklesparkle|t|0.2023|0.0|0.904|0.096|RT @MrBudSmith: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/8xo
AndrewR_Physics|ProfChrisMJones|0.0|0.0|1.0|0.0|"RT @ProfChrisMJones: As an academic, Trump's election was a wake-up call to me, but not for the reasons that @NickKristof seems to think. h"
tejana1234|summerbrennan|-0.4767|0.163|0.837|0.0|"RT @summerbrennan: As I've said before, I called McCain and Graham offices multiple times in tears right after the election and they are no"
BonnieGranny|hautedamn|-0.34|0.113|0.833|0.054|RT @hautedamn: The people who want you to believe Russia hacked the election are the same people telling you #pizzagate isn't real.
FrankDObrad|twitter|-0.25|0.1|0.9|0.0|I still find it a bit to coincidental that Hillary cancelled her fireworks display the day before the election. Som https://t.co/fldCv5NcDo
_dooooreen|vicenews|-0.3612|0.116|0.884|0.0|"RT @vicenews: I think its ridiculous"" Trump continues to shrug off a CIA report that Russia meddled in the 2016 election https://t.co/p6m"
_dooooreen|t|-0.3612|0.116|0.884|0.0|"RT @vicenews: I think its ridiculous"" Trump continues to shrug off a CIA report that Russia meddled in the 2016 election https://t.co/p6m"
AkaMotherto3|twitter|-0.2302|0.14|0.75|0.109|Sue to throw MI EC votes out. Or sue for hand count. This election is so screwed up. Include #putingate &amp; its tota https://t.co/iFI6PywAgn
christina_hikes|nytimes|0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
christina_hikes||0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
quailcrown|BrendanNyhan|-0.4659|0.169|0.787|0.043|"RT @BrendanNyhan: Seeing people dismiss as silly conspiracy talk, but far more serious. Potential Dep SOS suggesting Obama used IC in a dom"
Iam_Books|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
hheyitsmonica|HockeywthHannah|0.0|0.0|1.0|0.0|@HockeywthHannah shady: the theme of the election
manning1018|HaileeSteinfeld|0.6808|0.0|0.781|0.219|RT @HaileeSteinfeld: I choose to be optimistic &amp; hopeful regardless of the election results. Our future depends on us coming together &amp; fin
LoveShaneal|MarketWatch|0.5719|0.0|0.844|0.156|"RT @MarketWatch: There's one stock that was down 79% YTD before Trump won the election, and has rocketed 131% since: https://t.co/MRDTi3OA1c"
LoveShaneal|marketwatch|0.5719|0.0|0.844|0.156|"RT @MarketWatch: There's one stock that was down 79% YTD before Trump won the election, and has rocketed 131% since: https://t.co/MRDTi3OA1c"
GH_obsession|summerbrennan|-0.4767|0.163|0.837|0.0|"RT @summerbrennan: As I've said before, I called McCain and Graham offices multiple times in tears right after the election and they are no"
ChrisGaryL|MaxSteel747|-0.6908|0.231|0.769|0.0|RT @MaxSteel747: Democrats Are Using the Same Corrupt Political System to Steal the Presidency From Trump &amp; Claim Russians Rigged Election~
The_InMediasRes|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
BourneInTexas|NotJoshEarnest|-0.4738|0.206|0.702|0.092|"RT @NotJoshEarnest: Remember when not accepting election results was a danger to the democracy? Seems like it was last month. Oh wait, it w"
Woolndoghairs|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
Woolndoghairs||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
Anyshka|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
KevinGFox|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
MEMasciale|nytimes|0.4939|0.0|0.686|0.314|"Russias Hand in Americas Election, via @nytimes https://t.co/VpvuxTOtxF"
MEMasciale|nytimes|0.4939|0.0|0.686|0.314|"Russias Hand in Americas Election, via @nytimes https://t.co/VpvuxTOtxF"
CharlesHamerle|laurahollis61|-0.6486|0.238|0.762|0.0|"RT @laurahollis61: This whole ""Russians hacked the election"" story is the biggest load of crap since#Benghazi ""it-was-a-video."" Dems are d"
klormpster|_Makada_|-0.296|0.115|0.826|0.06|"RT @_Makada_: President-Elect Trump: It's ridiculous to say Russia intervened in the election, I think it's just another excuse. We had a m"
JoseyOhh|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
Glen_Coco2193|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
knowlton_paula|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
guna15|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
sumoh7|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
sumoh7|change|0.0|0.0|1.0|0.0|RT @starfirst: 2016 Presidential Election Results May be Invalid https://t.co/ZjJBAAj53J via @Change
InChargeable1|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
ElaineFox|SocialNews|0.0|0.0|1.0|0.0|RT @SocialNews: Russian 'Meddling' In Election: Most Overblown Story Ever? https://t.co/iOIb10ZL3L
ElaineFox|powerlineblog|0.0|0.0|1.0|0.0|RT @SocialNews: Russian 'Meddling' In Election: Most Overblown Story Ever? https://t.co/iOIb10ZL3L
Acliffe|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/DCotOqPic0 https://t."
Acliffe||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/DCotOqPic0 https://t."
SandiChilds|swin24|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
SandiChilds|thedailybeast|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
clausen_ed|politico|0.0|0.0|1.0|0.0|RT @politico: .@SenSchumer demands congressional inquiry on Russian meddling https://t.co/eD2nlokARd https://t.co/Uk7ShnuCEj
clausen_ed|politico|0.0|0.0|1.0|0.0|RT @politico: .@SenSchumer demands congressional inquiry on Russian meddling https://t.co/eD2nlokARd https://t.co/Uk7ShnuCEj
iNewsSource|DefenseOne|0.0|0.0|1.0|0.0|RT @DefenseOne: Obama Orders 10-Year Deep Dive into Election Hacking https://t.co/QIH0t8awqU | @DefTechPat https://t.co/66x7iYcz80
iNewsSource|defenseone|0.0|0.0|1.0|0.0|RT @DefenseOne: Obama Orders 10-Year Deep Dive into Election Hacking https://t.co/QIH0t8awqU | @DefTechPat https://t.co/66x7iYcz80
sponson|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
sponson|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
rickybobby90210|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
rickybobby90210|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
GraggQuinton|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
GraggQuinton|t|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
Paratisi|hautedamn|-0.34|0.113|0.833|0.054|RT @hautedamn: The people who want you to believe Russia hacked the election are the same people telling you #pizzagate isn't real.
mcormack1977|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
THAToneil|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
camper_bruce|hautedamn|-0.34|0.113|0.833|0.054|RT @hautedamn: The people who want you to believe Russia hacked the election are the same people telling you #pizzagate isn't real.
stevieboy13|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ShainEThomas|JuddLegum|-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
ShainEThomas||-0.5081|0.12|0.88|0.0|RT @JuddLegum: 3. He went on TV today with an absolutely insane theory: it wasn't Russia behind the election hacks -- it was Obama! https:/
neurotrade|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
britswitz|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
littleponies|YouTube|0.0|0.0|1.0|0.0|Eric Shawn reports: The alleged Russian election hacking https://t.co/uv7Xv0ms6V via @YouTube
littleponies|linkis|0.0|0.0|1.0|0.0|Eric Shawn reports: The alleged Russian election hacking https://t.co/uv7Xv0ms6V via @YouTube
ambersimmons26|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
NCPatriotMom|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
NCPatriotMom|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
ralphharper1965|ucbearcats1|0.0|0.0|1.0|0.0|"RT @ucbearcats1: @RBReich From the Emoluments clause to Russia hacking the election, #ComradeTrump is not properly qualified to be Presiden"
JBax52|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Peresson79|nanakim07|0.0|0.0|1.0|0.0|RT @nanakim07: https://t.co/qwjT0ZEzYH
Peresson79|cnn|0.0|0.0|1.0|0.0|RT @nanakim07: https://t.co/qwjT0ZEzYH
RussellSaylor|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
film_planet|Boofyre|-0.1027|0.11|0.8|0.09|RT @Boofyre: Police admit sex complaint against Assange was fabricated in elaborate plot https://t.co/O5quK6z26O ... by #ProgressiveShay vi
film_planet|linkis|-0.1027|0.11|0.8|0.09|RT @Boofyre: Police admit sex complaint against Assange was fabricated in elaborate plot https://t.co/O5quK6z26O ... by #ProgressiveShay vi
ZappaSzep|kjacobsedits|0.4574|0.0|0.85|0.15|RT @kjacobsedits: Looking for a pro-women organization you can support in the wake of the election? Try @girlswritenow! https://t.co/YyljR7
ZappaSzep|t|0.4574|0.0|0.85|0.15|RT @kjacobsedits: Looking for a pro-women organization you can support in the wake of the election? Try @girlswritenow! https://t.co/YyljR7
ellen_ritt|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
Zhian2160|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Other than @LindseyGrahamSC is there a single principled Republican in Washigton? Russia directly intervened in our electio
MelanieKV|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
KingisPingis|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
brandon_fields|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
pgrandee10|1fourallfour1|-0.1613|0.163|0.706|0.131|RT @1fourallfour1: This ain't over folks we WON'T accept RIGGED election #Resist #AuditTheVote #Recount2016 #TheResistance #notmypresident
vivs1man|rwindrem|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
vivs1man|nbcnews|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
KathleenELoughr|TeaPainUSA|-0.4215|0.141|0.859|0.0|"RT @TeaPainUSA: This is the first election in American history that the incoming President is the ""lame duck."""
ToddDomke|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
dell_cheryl|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
AndreFrato|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
AndreFrato|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
ElizbethLManess|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
hexogennotsugar|mhmck|0.0|0.0|1.0|0.0|"RT @mhmck: Rerun the election. Paper ballots. Two names: Clinton, Trump. International observers by the tens of thousands. Ukraine did it."
tptdave|emigre80|-0.3802|0.217|0.662|0.121|"RT @emigre80: Both Trump and Sanders were delighted to cry ""rigged election!"" when they ran against Clinton.Now that there's evidence? *C"
macvolley1|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
JJFan18|JuddLegum|0.4404|0.0|0.847|0.153|RT @JuddLegum: Updated list of GOP members supporting investigation into Russian interference w/prez electionSen GrahamSen McCainSen Co
USA_Jedi|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
EnarDavis1|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
FlorianM1_|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
wtflanksteak|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
poodbit499|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
CrystalEffect_|YouTube|-0.2342|0.242|0.614|0.143|I liked a @YouTube video from @jaclynglenn https://t.co/PWdyx0ismJ Girl FREAKS OUT over Donald Trump losing the election
CrystalEffect_|youtube|-0.2342|0.242|0.614|0.143|I liked a @YouTube video from @jaclynglenn https://t.co/PWdyx0ismJ Girl FREAKS OUT over Donald Trump losing the election
Paratisi|CourageOfWisdom|-0.6153|0.216|0.676|0.108|"RT @CourageOfWisdom: GRAHAM &amp; McCAIN, MOST CORRUPT &amp; EVIL SENATORS IN D.C. Gaslighting Americans is a HUGE misuse of power. #pizzagate http"
BenBergerBaby|vicenews|-0.3612|0.116|0.884|0.0|"RT @vicenews: I think its ridiculous"" Trump continues to shrug off a CIA report that Russia meddled in the 2016 election https://t.co/p6m"
BenBergerBaby|t|-0.3612|0.116|0.884|0.0|"RT @vicenews: I think its ridiculous"" Trump continues to shrug off a CIA report that Russia meddled in the 2016 election https://t.co/p6m"
PBG2017|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
PBG2017|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
Allnkat|washingtonpost|-0.2732|0.14|0.726|0.134|She is laughable:         Kellyanne Conway calls CIA report on Russian election meddling laughable and ridiculous https://t.co/q1ivm7KKxA
FlyingYogini|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
Serabbi|politicususa|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
Serabbi|twitter|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
xxdesmus|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
xxdesmus|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
MexicanCareBear|BardockObama|-0.8208|0.322|0.591|0.087|"RT @BardockObama: Liberals are so stupid y'all ask for a recount then fail, then think Russia rigged the election lol it was obviously J Co"
kentrmoore|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
MiamiDadeFLA|tkinder|-0.3182|0.134|0.802|0.064|RT @tkinder: Kellyanne Conway calls CIA report on Russian election meddling 'laughable and ridiculous' - https://t.co/p3hWPT87in via @nuzzel
MiamiDadeFLA|washingtonpost|-0.3182|0.134|0.802|0.064|RT @tkinder: Kellyanne Conway calls CIA report on Russian election meddling 'laughable and ridiculous' - https://t.co/p3hWPT87in via @nuzzel
tadpoledrain|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
TRAPCASH|SenatorTomUdall|0.5267|0.067|0.714|0.219|RT @SenatorTomUdall: I will join lawmakers in both parties &amp; demand investigation of Russia's effort to influence presidential election. ht
KTynot|DonaldJFunk|-0.1685|0.089|0.911|0.0|RT @DonaldJFunk: Incredible that Obama hasn't launched full investigation of Comey &amp; Russian interference w/ election! @ezlusztig @kurteich
tkdcoach|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
merryannmariano|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
merryannmariano|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
SOcean5|hale_razor|-0.4033|0.181|0.738|0.081|RT @hale_razor: Leftists very concerned Trump may be cozy with Russia had no problem with Obama telling Putin he'll be more flexible after
slickvolt|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
No_Kipling|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
No_Kipling|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
JanettePattison|EcuadorDeb|0.0|0.0|1.0|0.0|RT @EcuadorDeb: @Irwin_Elaine @_0HOUR1 Shows that if Putin really wanted to influence the election all he had to do was donate to the Clint
jjj5819|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Wjdiaz1965|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
575haiku|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
janinewallace|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
billm9|WSJ|0.0|0.0|1.0|0.0|Georgia reported an attempt to hack its election database via a U.S. government IP address  https://t.co/4rHQ7yMukQ via @WSJ
billm9|wsj|0.0|0.0|1.0|0.0|Georgia reported an attempt to hack its election database via a U.S. government IP address  https://t.co/4rHQ7yMukQ via @WSJ
mikegraham57|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
PressRevere|paulareverepress|0.0|0.0|1.0|0.0|Founding Fathers Say Russia Election Interference Means Electoral College Must RejectTrump https://t.co/N0aBE3RzRP https://t.co/6g2ZNcu8OT
srchadaga|SenatorTomUdall|0.5267|0.067|0.714|0.219|RT @SenatorTomUdall: I will join lawmakers in both parties &amp; demand investigation of Russia's effort to influence presidential election. ht
toussaintgroup|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
toussaintgroup||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
ellehilley|_discosuperfly_|0.3612|0.0|0.815|0.185|RT @_discosuperfly_: if only Michigan looked like this during the election https://t.co/VW1jckKlQD
ellehilley|twitter|0.3612|0.0|0.815|0.185|RT @_discosuperfly_: if only Michigan looked like this during the election https://t.co/VW1jckKlQD
JoyRedeemed|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
JoyRedeemed||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
deborahjlundy|ProgressiveShay|-0.7579|0.338|0.597|0.065|RT @ProgressiveShay: @kierobar THIS is scary as shit. They want to discredit the election. omg.
zeering_road|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
zeering_road|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
annendress|twitter|0.4404|0.0|0.847|0.153|I hope voter ID becomes the law so we don't have to go thru this next election https://t.co/NTUZwUnhgS
thejohnbondshow|EllenMeister|0.0|0.0|1.0|0.0|@EllenMeister Democrats have been importing foreign influence in our election process through mass immigration for 50 years.
srikki03|igorvolsky|-0.2732|0.123|0.877|0.0|RT @igorvolsky: Putting the GOP's complete disregard for Putin's meddling in our election into context. https://t.co/xgffbrjk81
srikki03|twitter|-0.2732|0.123|0.877|0.0|RT @igorvolsky: Putting the GOP's complete disregard for Putin's meddling in our election into context. https://t.co/xgffbrjk81
3045hobart|raymondjlee|0.4588|0.0|0.81|0.19|RT @raymondjlee: Dear @POTUS @SenateDems @HouseDemocrats If there's been evidence of election tampering can we finally legally take action
KoalaBerries|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
RobertLeydon|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
NancyDiMattia1|ErnestRickard|0.0|0.0|1.0|0.0|RT @ErnestRickard: Sign the petition to overturn the  #Overturn2016PresElection  https://t.co/fufOmPb8ir
NancyDiMattia1|petitions|0.0|0.0|1.0|0.0|RT @ErnestRickard: Sign the petition to overturn the  #Overturn2016PresElection  https://t.co/fufOmPb8ir
kcnewhaven|JohnWDean|0.0|0.0|1.0|0.0|RT @JohnWDean: The intel report on Russia's role in the 2016 election must be available for all electors before the electoral college meets
slidewinding|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
slidewinding|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
mjohnso27|ericgarland|0.0|0.0|1.0|0.0|RT @ericgarland: Do you tell America the day after the election that Russia spearfished all of our think tanks in brazen fashion?
wifflewaffel|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
wifflewaffel|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
annabelslil|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
EryckahAnne|ParkerMolloy|-0.5067|0.17|0.83|0.0|"RT @ParkerMolloy: ""patrioteagle.flag says there's a child sex pizza dungeon!""""On it!""""The CIA says Russia messed w/ the election!""Some s"
Hefflin|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
626__624|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
peruchin54|newcenturytimes|0.0|0.0|1.0|0.0|https://t.co/XkqRu5efXb
tardiskitten|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
JPReed92|thetrudz|-0.2263|0.122|0.751|0.127|"RT @thetrudz: Every time a cowardly White liberal writes a ""coddle bigots, already"" defense of White supremacy article post-election, my mi"
jordan_erdakos|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
anticorrup_coah|PrisonPlanet|-0.5106|0.191|0.809|0.0|"RT @PrisonPlanet: Post election riots: FAILED.Jill Stein recount: FAILED.Intimidation of EC members: FAILED.""Fake news"": FAILED.""Russia"
tarttwit|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
InvestInDenim|FieryRedReviews|0.6486|0.137|0.474|0.389|RT @FieryRedReviews: Please sign to help save our country from fascism and treason: https://t.co/vxhcIfe5Qp
InvestInDenim|petitions|0.6486|0.137|0.474|0.389|RT @FieryRedReviews: Please sign to help save our country from fascism and treason: https://t.co/vxhcIfe5Qp
JackMartin96763|NCbgirl|0.0|0.0|1.0|0.0|RT @NCbgirl: @MaydnUSA @LIpatriot1 - REMEMBER THIS?Talk about interfering in another country's election . . . https://t.co/VhofKRLLLM
JackMartin96763|twitter|0.0|0.0|1.0|0.0|RT @NCbgirl: @MaydnUSA @LIpatriot1 - REMEMBER THIS?Talk about interfering in another country's election . . . https://t.co/VhofKRLLLM
JuliaGS|MarkSimoneNY|-0.197|0.075|0.925|0.0|"RT @MarkSimoneNY: Hillary looks the other way when Russia invades countries, sells them 25% of our uranium. So they rig the election agains"
EzabQuader|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
Mo_An2016|HispanicsTrump|0.0|0.0|1.0|0.0|RT @HispanicsTrump: If Hillary really wants to know who cost her the election all she needs to do is look in the mirror... #FakeNews #Russi
dianemcaul|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Landwehr_Erik|GeorgeTakei|-0.4199|0.108|0.892|0.0|"RT @GeorgeTakei: Mitch McConnell tried to cast doubt on the CIA findings before the election. Then, magic! His wife Elaine Chao is named Tr"
tonecky|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
DJT_ChosenbyGod|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
DJT_ChosenbyGod|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
momof3moochers|foxnation|0.0|0.0|1.0|0.0|"RT @foxnation: .@JudgeJeanine: The Election Is Over, Mr. President https://t.co/VW0vBabMjz"
momof3moochers|nation|0.0|0.0|1.0|0.0|"RT @foxnation: .@JudgeJeanine: The Election Is Over, Mr. President https://t.co/VW0vBabMjz"
independentpen|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
BelewforSheriff|nbc29|0.7088|0.0|0.743|0.257|Good Evening! On January 10th there will be a special election to replace Tom Garrett in the Virginia State... https://t.co/o3zc1cmpcy
pmcall|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
pmcall|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
TYdal_wave7844|swin24|-0.0572|0.055|0.945|0.0|"RT @swin24: Today, Trump says he doesnt want anyone hacking the U.S.In July, he called on Russia to hack the U.S. govt.https://t.co/"
PaulaBuermele|TinyTinyTrump|0.5635|0.14|0.495|0.365|"@TinyTinyTrump @Bill_Rhodes54 Well, they weren't smart enough to win the election."
RRMGOP|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
BoxANT|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
BoxANT|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
JuliaR1414|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Iamnowblue|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
Iamnowblue||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
viptandon|slone|0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
viptandon||0.6714|0.0|0.8|0.2|RT @slone: GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.c
Alice16050204|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
TeamTrumpTeX|MissLizzyNJ|-0.952|0.53|0.47|0.0|"RT @MissLizzyNJ: #ImStillNotOver the fact that I lost the election because I'm a lying criminal and America hates me, so I'll blame fake ne"
runningwnails|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
cant_king|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
mchwllms5|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
SandiChilds|swin24|-0.0572|0.055|0.945|0.0|"RT @swin24: Today, Trump says he doesnt want anyone hacking the U.S.In July, he called on Russia to hack the U.S. govt.https://t.co/"
jalivezb|Phaedrus08|-0.6144|0.277|0.625|0.098|@Phaedrus08 @goodtroubleme @VABVOX @BernieSanders I don't remember him losing 2 a racist Cheeto n a gimme election. Then hiding in the woods
Atticus_Amber|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
NancyBess|Pinkcloud15|0.2225|0.0|0.914|0.086|RT @Pinkcloud15: It's time 2 take our country back! Call the W H 202-456-1414 'n tell thm U want a new election done w/paper ballots! https
LordDayoo|FoxNews|0.0|0.0|1.0|0.0|RT @FoxNews: U.S. markets since election. https://t.co/NRw2LedQ7u
LordDayoo|twitter|0.0|0.0|1.0|0.0|RT @FoxNews: U.S. markets since election. https://t.co/NRw2LedQ7u
JC12Tx|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
stgrizelda|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
mamalocaz|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
steph_bello|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
maketrumpgoaway|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
maketrumpgoaway|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
KnowledgIsPowa|aliasvaughn|-0.2263|0.087|0.913|0.0|RT @aliasvaughn: This petition demanding a new election with paper ballots needs 100k signatures before EC votes. If you can spare a minute
AustinTG_15|Kasper_Tait|0.2406|0.165|0.638|0.197|RT @Kasper_Tait: russia hey u hacked the election results could u maybe hack my bank account. . . like add a few more zeros or ?? haha no p
mrfusspot|mtracey|0.0|0.0|1.0|0.0|"@mtracey If they can prove the Russians did the election, can we just get a new set of candidates to vote for?"
mjohnso27|ericgarland|-0.296|0.099|0.901|0.0|RT @ericgarland: Do you come out the day after this totally weird-smelling abomination of an election with all its technical difficulties?
JPReed92|thetrudz|-0.0299|0.09|0.824|0.086|"RT @thetrudz: It is Whites who've ignored who we are, not the other way around. Don't let these cowardly White liberal post-election articl"
e_revolutionist|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
GL_Funky|dylanmarron|-0.3802|0.126|0.874|0.0|"RT @dylanmarron: Liberal Professor in @nytimes: ""Push for trans rights lost us the election!""Reality: Anti-trans bathroom laws make N.C."
momof3moochers|FoxNews|0.1027|0.089|0.806|0.105|"RT @FoxNews: Last night on ""Justice,"" @JudgeJeanine had stark words for those who refuse to accept the results of the election. https://t.c"
momof3moochers||0.1027|0.089|0.806|0.105|"RT @FoxNews: Last night on ""Justice,"" @JudgeJeanine had stark words for those who refuse to accept the results of the election. https://t.c"
Sparblack1213|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
Sparblack1213|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
vivigold197|MrDane1982|-0.3716|0.139|0.861|0.0|RT @MrDane1982: Bernie Sanders and Donald Trump were both screaming the election was rigged but now Bernie is mute and Trump is in denial a
clausen_ed|swin24|0.6369|0.0|0.755|0.245|"RT @swin24: Trump '12/'14: bashes Obama 4 skipping intel briefingsTrump now: I skip briefings cuz Im, like, a smart person https://t.c"
clausen_ed||0.6369|0.0|0.755|0.245|"RT @swin24: Trump '12/'14: bashes Obama 4 skipping intel briefingsTrump now: I skip briefings cuz Im, like, a smart person https://t.c"
calRINOhunter|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
rhondastew|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
Teri_A_Adams|tamisflo65|-0.5267|0.139|0.861|0.0|"RT @tamisflo65: @VictorB123 @Ktrotter80 Victor, it's not about the election. It's about a threat to our country. Do you not see that? @Lane"
JustMeinMI|twitter|0.4877|0.0|0.851|0.149|"So many Trump supporters assumed he'd become presidential after the election. This is as presidential as it gets, a https://t.co/rlkKfFyeBK"
tealalltheway|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
tealalltheway|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
antiqueseahorse|NinjaEconomics|0.0|0.0|1.0|0.0|"RT @NinjaEconomics: NPR has independently confirmed the CIA's new assessment that ""Russia was trying to tip the election to Trump."" https:/"
antiqueseahorse||0.0|0.0|1.0|0.0|"RT @NinjaEconomics: NPR has independently confirmed the CIA's new assessment that ""Russia was trying to tip the election to Trump."" https:/"
ZalMox3|Kasparov63|0.2263|0.0|0.899|0.101|RT @Kasparov63: I wrote many columns about Trump &amp; Putin's involvement in the election all year. Worth revisiting. https://t.co/IFEFu6SaMk
ZalMox3|huffingtonpost|0.2263|0.0|0.899|0.101|RT @Kasparov63: I wrote many columns about Trump &amp; Putin's involvement in the election all year. Worth revisiting. https://t.co/IFEFu6SaMk
edgary1|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
rescuedogsrok|riotwomennn|0.296|0.0|0.879|0.121|"RT @riotwomennn: Russian Deputy Foreign Minister Sergei Ryabkov admits Russian gov ""maintained contacts"" w Trump during election  https://t"
rescuedogsrok||0.296|0.0|0.879|0.121|"RT @riotwomennn: Russian Deputy Foreign Minister Sergei Ryabkov admits Russian gov ""maintained contacts"" w Trump during election  https://t"
Jpdavi4|voxdotcom|0.0|0.0|1.0|0.0|"Russia's role in this year's presidential election, explained by a media historian https://t.co/jFBferyYZG via @voxdotcom"
Jpdavi4|vox|0.0|0.0|1.0|0.0|"Russia's role in this year's presidential election, explained by a media historian https://t.co/jFBferyYZG via @voxdotcom"
ABCVeterans2015|DeSmogCanada|0.0|0.0|1.0|0.0|RT @DeSmogCanada: I dont think they wanted to kick us out during the election campaign. https://t.co/NrU6EB8vNa #bcpoli #cdnpoli #SiteC
ABCVeterans2015|desmog|0.0|0.0|1.0|0.0|RT @DeSmogCanada: I dont think they wanted to kick us out during the election campaign. https://t.co/NrU6EB8vNa #bcpoli #cdnpoli #SiteC
nw_deplorable|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
billm9|veggie64_leslie|-0.3016|0.145|0.759|0.096|"RT @veggie64_leslie: Homeland Security IP address linked to attempted hack into GA voting systemIs this ""fake news"" HRC was afraid of?htt"
MattyPGood|leahmcelrath|0.5584|0.0|0.796|0.204|RT @leahmcelrath: Watergate seems like such an minor almost innocent bit of subterfuge compared to what's happened in this election.
Elizabeth_J91|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
chaquewe7|politico|0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
chaquewe7||0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
Scout2462|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
wonggal|twitter|0.3612|0.0|0.8|0.2|seems like every day produces another irregularity about prez election....sigh... https://t.co/4F0QAz7M4Y
eddie736|okrent|0.0|0.0|1.0|0.0|"RT @okrent: Trump transition team: ""The election ended...in one of the biggest Electoral College victories in history."" Right - 46th larges"
zunderwhelmed|bravenew1|0.5859|0.0|0.798|0.202|"RT @bravenew1: FBI covered up Russian influence on Trump's election win, Harry Reid claims https://t.co/KmdByXfok4 #InvalidElection"
zunderwhelmed|theguardian|0.5859|0.0|0.798|0.202|"RT @bravenew1: FBI covered up Russian influence on Trump's election win, Harry Reid claims https://t.co/KmdByXfok4 #InvalidElection"
StoneColdChik|StoneColdChik|-0.4939|0.158|0.842|0.0|RT @StoneColdChik: this is hillary obama mccain graham burr and this administration attempting to steal the election https://t.co/FsC7FQ1FEG
StoneColdChik|rt|-0.4939|0.158|0.842|0.0|RT @StoneColdChik: this is hillary obama mccain graham burr and this administration attempting to steal the election https://t.co/FsC7FQ1FEG
r1965rainey|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
kemalkirisci|BrookingsInst|0.0|0.0|1.0|0.0|RT @BrookingsInst: 46% of Americans think Obama should take action on Israel-Palestine before leaving office https://t.co/pr01irnpBj https:
kemalkirisci|brookings|0.0|0.0|1.0|0.0|RT @BrookingsInst: 46% of Americans think Obama should take action on Israel-Palestine before leaving office https://t.co/pr01irnpBj https:
AllDayAMazing|timcarvell|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
AllDayAMazing|freep|-0.1531|0.143|0.738|0.119|RT @timcarvell: @markoff 4. The actual situation is bad enough w/o needing to hype it up. Better article here: https://t.co/QKF8lsoHJw
Gary_Davis_7807|abermans|-0.3802|0.126|0.874|0.0|RT @abermans: 2/2017 #Election?Come what #may wants:More #Brexit delay and more tory power.Only she will get mass #UKIP upvote!https://
Gary_Davis_7807||-0.3802|0.126|0.874|0.0|RT @abermans: 2/2017 #Election?Come what #may wants:More #Brexit delay and more tory power.Only she will get mass #UKIP upvote!https://
jrrom|laurahollis61|-0.6486|0.238|0.762|0.0|"RT @laurahollis61: This whole ""Russians hacked the election"" story is the biggest load of crap since#Benghazi ""it-was-a-video."" Dems are d"
JJFan18|jkarsh|0.4576|0.0|0.87|0.13|"RT @jkarsh: Given the CIA report about Russia influencing our election, this line from an @azcentral piece is very interesting. https://t.c"
JJFan18||0.4576|0.0|0.87|0.13|"RT @jkarsh: Given the CIA report about Russia influencing our election, this line from an @azcentral piece is very interesting. https://t.c"
HahnAmerica|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
gurusix|pattonoswalt|0.4939|0.0|0.882|0.118|"RT @pattonoswalt: Seems to me, you didn't wanna talk about it before the election. Seems to me, you just turned your pretty head &amp; walked a"
StarCityBFFs|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
A_HolePatrol|pattonoswalt|0.4939|0.0|0.882|0.118|"RT @pattonoswalt: Seems to me, you didn't wanna talk about it before the election. Seems to me, you just turned your pretty head &amp; walked a"
CindyMae65|LindaSuhler|-0.2168|0.144|0.75|0.106|RT @LindaSuhler: Remember Obama's hot mic msg to Putin about flexibility after the election?What are they scared of? #RussianHackinghttps
crosa1988|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: BREAKING: Harry Reid says FBI Director James Comey deliberately withheld info on Russia's election meddling &amp; should re
PeabsLord|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: @EBrooksUncut Constitution. When election thrown into the House, the House elects the president. Can be anybody. For th"
rich_norseman22|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
glajchs|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
PiratesWife82|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
npnikk|npnikk|-0.5904|0.168|0.832|0.0|"RT @npnikk: Trump bashes CIA, dismisses Russian hacking report = FAKE NEWS -&gt; CIA cannot operate inside USA 2 produce report.. https://t.co"
npnikk|t|-0.5904|0.168|0.832|0.0|"RT @npnikk: Trump bashes CIA, dismisses Russian hacking report = FAKE NEWS -&gt; CIA cannot operate inside USA 2 produce report.. https://t.co"
pinkmartini12|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
geraldpayne25|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
lordsutch|trumwill|-0.1027|0.057|0.943|0.0|"RT @trumwill: If the election had been held  on that day, turnout would have been hard to gage because nobody would have known. https://t.c"
lordsutch||-0.1027|0.057|0.943|0.0|"RT @trumwill: If the election had been held  on that day, turnout would have been hard to gage because nobody would have known. https://t.c"
Zenkitty714|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
periodicaI|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/uRPI8WAryY
emccoy_writer|markberman|0.0|0.0|1.0|0.0|"RT @markberman: President-elect Trump, speaking to Fox News yesterday, again says he doesn't think Russia meddled in the election/doesn't t"
UserGlobal|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/7mF7q1Juo0
Amit258Rai|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
BostonDaveOH|RepublicanChick|-0.1779|0.082|0.918|0.0|"RT @RepublicanChick: Liberals are accusing Russia of influencing the election. At the same time, liberals enabled citizens of other countri"
NTrexit|Khanoisseur|0.5106|0.0|0.845|0.155|RT @Khanoisseur: .@LindseyGrahamSC Strong bipartisan statement on Russian meddling in election But you all need to also investigate FBI i
starrhaus|scottwongDC|-0.34|0.112|0.888|0.0|"RT @scottwongDC: In rare bipartisan statement, McCAIN, GRAHAM, SCHUMER &amp; REED say reports of Russian interference in election ""should alarm"
mekmtl|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
sylviapataki|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
designergrace|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
Oliver_Zhang_|Holbornlolz|-0.6705|0.231|0.684|0.085|RT @Holbornlolz: People who killed 100's of 1000's to ensure regime change all over the M. East are upset that Russia may have interfered i
bstrand|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
bstrand|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
butte_tocks|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
butte_tocks||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
terebifunhouse|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
terebifunhouse|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
hi_hat_truth|theonlyadult|0.0|0.0|1.0|0.0|@theonlyadult @nytimes why are the election results still being considered valid?
mortermermouse|chriscoxcountry|0.0|0.0|1.0|0.0|RT @chriscoxcountry: WeAll SHOULD BeAngry #VERYangry Bipartisan+anger+grows+over+Russian+interference+into+U.S.+election https://t.co/EMmjE
mortermermouse|t|0.0|0.0|1.0|0.0|RT @chriscoxcountry: WeAll SHOULD BeAngry #VERYangry Bipartisan+anger+grows+over+Russian+interference+into+U.S.+election https://t.co/EMmjE
1Luv2|leahmcelrath|-0.3412|0.112|0.888|0.0|RT @leahmcelrath: NYTimes Editorial Board takes a stand &amp; even calls Trump out for not supporting an investigation into Russia hackinghttp
sasyecat|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
FairmanAngel|AnnaSophia_TOPS|-0.8264|0.278|0.722|0.0|RT @AnnaSophia_TOPS: Wasn't it some dems that hacked the election w/all their CHEATING? What about that? 50+ yrs too! Project Veritas vids
MadJewessWoman|MadJewessWoman|0.0|0.0|1.0|0.0|"RT @MadJewessWoman: .@realDonaldTrumpINVESTIGATE @SenJohnMcCain 4 overthrowing #Ukraine govt, influencing election in #KIEV, 2013-14http"
CVoelkerding|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
linksteroh|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
linksteroh||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
slone|realDonaldTrump!!!|0.6714|0.0|0.78|0.22|GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.co/uteNKYRWWo
slone|nbcnews|0.6714|0.0|0.78|0.22|GOOD CHOICE @realDonaldTrump!!! Rex Tillerson of ExxonMobil Expected to Be Named Trump's Secretary of State: Sources https://t.co/uteNKYRWWo
dbergg|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
dbergg|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
BellTrumpkin|carolinagirl217|-0.6808|0.397|0.603|0.0|RT @carolinagirl217: Outrageous:-Debt-Benghazi-ACA-Increased Terrorism -Emails-Iran-Govt Overreach/EO-Riots-Fake MSM Newshttps:
JeromeDawson3|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
JeromeDawson3|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
jmlara02|LeahR77|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
jmlara02|t|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
DockedinNewYork|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
MissKittyfromVa|laurahollis61|-0.6486|0.238|0.762|0.0|"RT @laurahollis61: This whole ""Russians hacked the election"" story is the biggest load of crap since#Benghazi ""it-was-a-video."" Dems are d"
Holmesdonna1|charliekirk11|-0.7184|0.269|0.731|0.0|RT @charliekirk11: Democrats blame the Russians and the FBI for their election loss. Was is the Russians that ignored middle America for
JackIrvin_RVA|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
JackIrvin_RVA||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
JoanieChesnutt|EcuadorDeb|0.0|0.0|1.0|0.0|RT @EcuadorDeb: @Irwin_Elaine @_0HOUR1 Shows that if Putin really wanted to influence the election all he had to do was donate to the Clint
bitznews|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/fyPkWvuKv0
reasonandlogic|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
AnnBGelder|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
SecurityKit|securitykit|-0.296|0.155|0.845|0.0|Obama orders review of election hacks as Trump doubts Russias role https://t.co/POuH4hCJ2A  #security
VinylQueen84|michaelianblack|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
VinylQueen84|twitter|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
konrad_jeff|JuddLegum|0.0|0.0|1.0|0.0|RT @JuddLegum: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/oRUPSkz7NV https:
konrad_jeff|medium|0.0|0.0|1.0|0.0|RT @JuddLegum: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/oRUPSkz7NV https:
NDgradmom|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
mr_boeb|jahimes|0.6375|0.0|0.754|0.246|RT @jahimes: @GoodJobGuru @PoliticalLine Yes. The election is over. But the electoral college has not met. So no President has been legally
clark7950|tteegar|-0.5242|0.232|0.67|0.098|RT @tteegar: BREAKING #RussianHackers made Hillary screech like an old crabby grandma &amp; lose the election!Nobody should be fooled! #Fak
SLadreda|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
SistaSoljaCtizn|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
bettyonline011|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
PubliusNV|MaryfromMarin|0.1007|0.125|0.729|0.145|RT @MaryfromMarin: @PubliusNV @WestDeclines Blame Melania! And Get Ready for the 'Post Trump' Haircut https://t.co/6BfncuqLSF #Election v
PubliusNV|pjmedia|0.1007|0.125|0.729|0.145|RT @MaryfromMarin: @PubliusNV @WestDeclines Blame Melania! And Get Ready for the 'Post Trump' Haircut https://t.co/6BfncuqLSF #Election v
DYoffee|LampOlive|-0.8004|0.255|0.745|0.0|RT @LampOlive: We all knew Trump couldn't win without rigging the election. Getting Russia to do it is the worst Avenue to go.
smokescreek|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
MarieMurcelle1|TomthunkitsMind|0.0|0.0|1.0|0.0|RT @TomthunkitsMind: Russia Says It Was In Touch With Trump Campaign During The Election. https://t.co/ik0yyqk7fF https://t.co/g7PF8uOlfg
MarieMurcelle1|huffingtonpost|0.0|0.0|1.0|0.0|RT @TomthunkitsMind: Russia Says It Was In Touch With Trump Campaign During The Election. https://t.co/ik0yyqk7fF https://t.co/g7PF8uOlfg
1finekitty|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
HonorFounders|HuffPostPol|-0.5719|0.252|0.748|0.0|Bipartisan anger grows over Russian interference into U.S. election https://t.co/325xuwbSHt via @HuffPostPol
HonorFounders|huffingtonpost|-0.5719|0.252|0.748|0.0|Bipartisan anger grows over Russian interference into U.S. election https://t.co/325xuwbSHt via @HuffPostPol
aringelestein|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
leoluminary|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
marymac169|ChicagoMGD|0.4767|0.0|0.853|0.147|RT @ChicagoMGD: @aliasvaughn @ezlusztig Reminder it isn't just the @CIA 16 other intelligence agencies had evidence of Russia's interferenc
vasilidante|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
vasilidante|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
madamecain|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
madamecain||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
Karenpacynski1|An0nKn0wledge|-0.6739|0.171|0.829|0.0|RT @An0nKn0wledge: THERE IS MORE EVIDENCE OF ALIENS EXISTING THEN THE RUSSIANS HACKING THE ELECTION.. BTW THE ELECTION FRAUD SO FAR ALL IN
hamel1776|youtube|0.0|0.0|1.0|0.0|CIA Splinter Group Calls For Overthrow Of Trump Election https://t.co/Kaazv6MvcI #YouTube #TheAlexJonesChannel
Landwehr_Erik|conlimonisal|0.0|0.0|1.0|0.0|"RT @conlimonisal: @Greg_Palast I don't understand why Hillary hasn't requested recount,considering all of the election tampering allegation"
SandiChilds|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
Changeisonus1|tonyschwartz|-0.4019|0.188|0.812|0.0|@tonyschwartz @1Luv2 An investigation is no substitute for a new election. The process was tainted and we demand a do-over.
TYdal_wave7844|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
snappyseaturtle|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
dindunuffinyt|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
dindunuffinyt|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
575haiku|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
575haiku|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
TynnaDemellier|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
alicia_bert|politicususa|0.4019|0.0|0.863|0.137|Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/Rf6JLQVQ9U
alicia_bert|politicususa|0.4019|0.0|0.863|0.137|Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/Rf6JLQVQ9U
mercedesfduran|bonita_jay1|0.0|0.0|1.0|0.0|"RT @bonita_jay1: @mercedesfduran @PattiKimble @JoyAnnReid I'm all for  that 1st choiceIn fact, here's a petition for another electn  https"
drmojo1975|LindaSuhler|-0.5574|0.247|0.753|0.0|RT @LindaSuhler: #FakeNews: CNN Shamed into Major Corrections on Ghana Election Storyhttps://t.co/czJezq4MlR
minirey805|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
minirey805|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
StevenChafin|ReveilleSoul1|-0.4019|0.119|0.881|0.0|"RT @ReveilleSoul1: This ""woman"" sets up a private server, aides running around w blackberrys full of state secrets &amp; cries Russia to overth"
THEJOKER20161|t|-0.3612|0.152|0.848|0.0|SKY SCUM VIEWS Trump: CIA Russia influence ridiculous https://t.co/kc6cR0ViSXIs the CIA investigating U2Knight of https://t.co/kRPg4KEu83
enolarae|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
enolarae||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Benjamin_T|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
The_ehrbaherba|thetrudz|-0.2263|0.122|0.751|0.127|"RT @thetrudz: Every time a cowardly White liberal writes a ""coddle bigots, already"" defense of White supremacy article post-election, my mi"
LyndasBags4fun|nytimes|0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
LyndasBags4fun||0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
caveboyjones|France4Hillary|0.0|0.0|1.0|0.0|RT @France4Hillary: BREAKING: Harry Reid says FBI Director James Comey deliberately withheld info on Russia's election meddling &amp; should re
bonniemac52|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
UnknownExtremes|mikeyymike78|0.0|0.0|1.0|0.0|RT @mikeyymike78: Major week in American politics coming up: Sec of State to be announced amid furor over reports Russia attempted to aide
juniperbreeze07|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
Annealeeb|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
suemagic|drjelks|-0.25|0.136|0.777|0.087|RT @drjelks: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/lGR9DEfPCL via @PalmerR
suemagic|palmerreport|-0.25|0.136|0.777|0.087|RT @drjelks: Michigan officials admit majority of Detroit vote counting machines broke on Election Day https://t.co/lGR9DEfPCL via @PalmerR
dr_tialynn|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
dr_tialynn||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
vivigold197|GareBearEsq|0.0|0.0|1.0|0.0|RT @GareBearEsq: Read this thread. And kunderstand that there are intel agents who know exactly what happened with our election. I said thi
pjmcgovern4|Watertowerjoey|-0.5267|0.216|0.784|0.0|"RT @Watertowerjoey: @kurteichenwald @rickitycrickety @infotrump2020 No, but the implication is that it turned the election.  No proof, yet"
freespeak3|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
pugewok|PowerPost|0.0|0.0|1.0|0.0|"RT @PowerPost: Key GOP senators call for bipartisan #Russia election probe, even as their leaders remain mum https://t.co/UOQqwDkbtN @elise"
pugewok|washingtonpost|0.0|0.0|1.0|0.0|"RT @PowerPost: Key GOP senators call for bipartisan #Russia election probe, even as their leaders remain mum https://t.co/UOQqwDkbtN @elise"
UppercutSlut|twitter|0.0772|0.112|0.762|0.126|"If anyone rigged the election it was Dems, not Russia. Trump should have had the popular vote too https://t.co/1Ka9nIKXA1"
304TheRevTJ|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
Destinyuhva|JoyAnnReid|0.4404|0.0|0.873|0.127|"RT @JoyAnnReid: Baer makes a good point: if we had been caught interfering in a foreign country's election, they would redo their election."
motatzin|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Kaladious|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
Kaladious|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
WayneSisk1|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
WayneSisk1||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
sumbodysbabygrl|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
dougnot2|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
dougnot2|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
yourbodybible|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
GreekSTL|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
PBPLife|theamericanmirror|0.0|0.0|1.0|0.0|Art of the deal... https://t.co/y7J4JPa2JN
NCPatriotMom|CDoranHarader|0.0|0.0|1.0|0.0|RT @CDoranHarader: CNN: Obama orders report into WikiLeaks timed for release just prior to Trump presidency https://t.co/pJZLWkJiWV ht... b
NCPatriotMom|linkis|0.0|0.0|1.0|0.0|RT @CDoranHarader: CNN: Obama orders report into WikiLeaks timed for release just prior to Trump presidency https://t.co/pJZLWkJiWV ht... b
metamemette|sethmoulton|0.6808|0.0|0.811|0.189|"RT @sethmoulton: Proud to see so many #MA6 constituents ready to work for change. There is so much to do, and this election was a call to a"
csittenfeld|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
csittenfeld|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
ENachmany|GovMikeHuckabee|0.3182|0.0|0.827|0.173|@GovMikeHuckabee Please the democrats will say anything to turn this election around
boandsunny|casatino|-0.1027|0.097|0.903|0.0|RT @casatino: FBI: sends vague letter; actually nothingMSM: *quivers*CIA: confirms Russia interfered w/electionMSM: \_()_/https://
cj15044|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
cj15044|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
aprov2480|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
aprov2480|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
K1er|tkinder|-0.3182|0.134|0.802|0.064|RT @tkinder: Kellyanne Conway calls CIA report on Russian election meddling 'laughable and ridiculous' - https://t.co/p3hWPT87in via @nuzzel
K1er|washingtonpost|-0.3182|0.134|0.802|0.064|RT @tkinder: Kellyanne Conway calls CIA report on Russian election meddling 'laughable and ridiculous' - https://t.co/p3hWPT87in via @nuzzel
kmclc2016brutus|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
suzykq5|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
JamesDubhthaigh|TheDailyEdge|-0.128|0.202|0.658|0.14|"RT @TheDailyEdge: RYAN (JUNE): ""We must stop cyber-attacks &amp; deliver justice to cyber assailants""CIA (DEC): Russia hacked the electionR"
GollyMollyB|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
ripple2012|cnn|0.0|0.0|1.0|0.0|Ex-CIA operative: We may need a new vote https://t.co/7JpmhboS9X
jglow70|SarahPalinUSA|-0.0422|0.118|0.77|0.112|RT @SarahPalinUSA: Russia's getting out of hand? So says the defeated. Not to worry... remember I can keep an eye on them from here. https:
NoveleraSalvaje|GeorgeTakei|0.0|0.0|1.0|0.0|"RT @GeorgeTakei: The CIA assessment concludes that Russians interfered with our election. With the margin so close, the result is illegitim"
wrdybrd|igorvolsky|-0.2732|0.123|0.877|0.0|RT @igorvolsky: Putting the GOP's complete disregard for Putin's meddling in our election into context. https://t.co/xgffbrjk81
wrdybrd|twitter|-0.2732|0.123|0.877|0.0|RT @igorvolsky: Putting the GOP's complete disregard for Putin's meddling in our election into context. https://t.co/xgffbrjk81
EnvyMeGreatly|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
leehlawrence|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/hMTCIFhYsd https://t."
leehlawrence||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/hMTCIFhYsd https://t."
zakbutterfield|rgodfrey|-0.0622|0.14|0.694|0.165|@rgodfrey I was so depressed after the election I forgot to thank you for serving the public on E-day. So I'm doing that now. Thank you.
cdelbrocco|m|-0.6342|0.207|0.793|0.0|He's a fucking liar!! Trump: It's 'Ridiculous' To Think Russia Intervened In The Election On My Behalf  https://t.co/hI0Wbo0CSd
molly_enselein|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
AnaCosentino2|dissentingj|0.296|0.178|0.593|0.229|@dissentingj @LyndaPole @CNBC @NBCNews No patience 4 Millennials..your protest vote handed election 2 Bozo.I hope you still like the circus
donna_king8|LibertyFolders|-0.5267|0.167|0.833|0.0|RT @LibertyFolders: Remember: Obama the hypocrite interfered in Israel's elections but he has balls 2 criticize Russia 4 supposedly interfe
davyd18|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
pinkmartini12|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
EffieGibbons|Lazarus1940|-0.34|0.13|0.87|0.0|"RT @Lazarus1940: @Sensiblecanadi1 @EffieGibbons @TheRebelTV @ibroxxxx @ezralevant CBC reported extensively on ""lake of fire"" comment in AB"
mjminpgh|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
lyoshki|SenatorTomUdall|0.5267|0.067|0.714|0.219|RT @SenatorTomUdall: I will join lawmakers in both parties &amp; demand investigation of Russia's effort to influence presidential election. ht
bachic2|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
biggsTRiPPYmane|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
2dJazz|koichinko|0.4588|0.0|0.833|0.167|Arc System Works Awards 2016 election results:GG: @koichinko &amp; @gou4th_fab BB: @soujif91 &amp; @MINAMI_IZANAMI Congr https://t.co/ywgd6kl4W6
2dJazz|twitter|0.4588|0.0|0.833|0.167|Arc System Works Awards 2016 election results:GG: @koichinko &amp; @gou4th_fab BB: @soujif91 &amp; @MINAMI_IZANAMI Congr https://t.co/ywgd6kl4W6
MtRushmore2016|NCbgirl|0.0|0.0|1.0|0.0|RT @NCbgirl: @MaydnUSA @LIpatriot1 - REMEMBER THIS?Talk about interfering in another country's election . . . https://t.co/VhofKRLLLM
MtRushmore2016|twitter|0.0|0.0|1.0|0.0|RT @NCbgirl: @MaydnUSA @LIpatriot1 - REMEMBER THIS?Talk about interfering in another country's election . . . https://t.co/VhofKRLLLM
afraud|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
SandiChilds|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
jwix57|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
PiratesWife82|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
PiratesWife82|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
LibertyBelle_76|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
dalydes|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
emzorbit|Bencjacobs|0.0|0.0|1.0|0.0|@Bencjacobs @pwthornton Casting shade. He has lit the fuse. Now any investigation into the election or DJT will erupt into a firestorm.
sasha031|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
sasha031|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
carlyandjack|twitter|-0.3147|0.222|0.778|0.0|Seriously! So now Obama sabotaged the election? Yikes! https://t.co/ILop2FVEHf
getrealvonciel|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
zeroinscw|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
zeroinscw|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
LukasZprehn|twitter|0.0|0.0|1.0|0.0|This is news to these people!? People who use the internet has known this since the first day of the election! Come https://t.co/vD3mtf5XFu
EmbryonicAttny|BryanDawsonUSA|-0.3612|0.135|0.865|0.0|RT @BryanDawsonUSA: GOP Congress:Hearings on #Benghazi witch hunt: 33Hearings on real Russian interference in US election: 0#russianha
realetybytes|Snap_Politics|0.0|0.0|1.0|0.0|RT @Snap_Politics: Speaking of foreign influences trying to throw US election.https://t.co/RpNwd85MCy#PaidBeatDowns at Trump rallies +Ele
janelleholmes20|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/4TnN8g6MGt https://t."
janelleholmes20||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/4TnN8g6MGt https://t."
marimegias|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
tifmcclure|DailyCaller|-0.6124|0.306|0.563|0.13|RT @DailyCaller: BuzzFeed Caught Citing Fake Data In Its Fake News Won The Election For Trump Argument  AGAIN https://t.co/5XVj30tggj ht
tifmcclure|dailycaller|-0.6124|0.306|0.563|0.13|RT @DailyCaller: BuzzFeed Caught Citing Fake Data In Its Fake News Won The Election For Trump Argument  AGAIN https://t.co/5XVj30tggj ht
NonCrystal|DanSlott|0.6124|0.0|0.783|0.217|RT @DanSlott: Imagine a thriller where at the climaxthe hero broadcasts a tape to the worldPROVING Russia fixed the U.S. election&amp; every
DirectorOfTech|mashable|0.0|0.0|1.0|0.0|RT @mashable: The one social platform actually taking action ahead of Trump's America https://t.co/4Q3d2SnM5G https://t.co/41TlUUVzx2
DirectorOfTech|mashable|0.0|0.0|1.0|0.0|RT @mashable: The one social platform actually taking action ahead of Trump's America https://t.co/4Q3d2SnM5G https://t.co/41TlUUVzx2
abbokey|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
luanph0311|MrBudSmith|0.2023|0.0|0.904|0.096|RT @MrBudSmith: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/8xo
luanph0311|t|0.2023|0.0|0.904|0.096|RT @MrBudSmith: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/8xo
blawgs_io|electionlawblog|-0.0772|0.098|0.902|0.0|Sorry But Alleged Russian Influence in Presidential Election Wont Lead to a Do-Over : https://t.co/MHsYqL0u3Y
mollymoor|BigRadMachine|0.5859|0.0|0.774|0.226|RT @BigRadMachine: The real winner of the election is every company that makes antidepressants.
soozanderson4|AG_Conservative|0.6124|0.115|0.577|0.308|RT @AG_Conservative: Both true:Russia actively worked to help Trump throughout election.HRC was an awful candidate who put own interest
soldierDtruth|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
deerhunter635|GitRDoneLarry|0.7084|0.124|0.612|0.264|RT @GitRDoneLarry: I know I said I'm blocking all Whiney election tweet but some are so dad gum entertaining! Ok starting again... now.
katherineislay|nytimes|0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
katherineislay||0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
McLonergan|LeahR77|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
McLonergan|t|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
Atheist_IMAGINE|kurteichenwald|-0.2382|0.22|0.67|0.11|"RT @kurteichenwald: No offense, @chucktodd, but when u say no one was sure Russia behind hack pre-election, shows u need to read more. http"
HostileParadox|EJDionne|0.0|0.0|1.0|0.0|"RT @EJDionne: ""Russia set out to influence the U.S. election..Republicans in Congress decided not to speak out against them..both calculati"
FelassanMa_lath|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
FelassanMa_lath|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Diannarinratmom|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
KweenLiapold|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
joanofarc1412|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
joanofarc1412|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
MtRushmore2016|LIpatriot1|0.5063|0.105|0.62|0.274|RT @LIpatriot1: @NCbgirl @MaydnUSA and if I'm not mistaken Obama played a hand in Canadian election
mellowkelo|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
mellowkelo||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
Ombudsman|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
BevPerryMusic|ProudlyLiberal2|0.0|0.0|1.0|0.0|"RT @ProudlyLiberal2: KeithOlbermann: This was not an election, this was a Coup D'Etat abetted by traitors. From 11/1: The Trumpchurian  ht"
birdsnfrogs|austinhollenba|-0.4215|0.141|0.859|0.0|"RT @austinhollenba: Here's the piece from the Detroit News, saying ""87 optical scanners broke on Election Day"" https://t.co/hGcHH5JN1v"
birdsnfrogs|detroitnews|-0.4215|0.141|0.859|0.0|"RT @austinhollenba: Here's the piece from the Detroit News, saying ""87 optical scanners broke on Election Day"" https://t.co/hGcHH5JN1v"
Twisty58|carold501|0.7881|0.143|0.515|0.342|"RT @carold501: Funny how the left laughed and said the election couldn't be hacked and then when their darling Hillary lost, they scream it"
clellab1|NotJoshEarnest|0.471|0.0|0.861|0.139|"RT @NotJoshEarnest: Listen up folks! Just because we lie about everything, doesn't mean we're lying about Russia hacking the election."
stldesktop|veggie64_leslie|-0.3016|0.145|0.759|0.096|"RT @veggie64_leslie: Homeland Security IP address linked to attempted hack into GA voting systemIs this ""fake news"" HRC was afraid of?htt"
alimhaider|Panhandlebound|0.0|0.0|1.0|0.0|@Panhandlebound EC either needs to overturn the election or we must redo the election https://t.co/eOpmTZ1mzt
alimhaider|cnn|0.0|0.0|1.0|0.0|@Panhandlebound EC either needs to overturn the election or we must redo the election https://t.co/eOpmTZ1mzt
SabrinaTenney|lindaantonO|0.0|0.0|1.0|0.0|@lindaantonO @Kriscental This is NOT about Hilary it's about another country hijacking our election.
herblatino|sunbeltgirl|-0.6478|0.202|0.798|0.0|"RT @sunbeltgirl: MT @INTJutsu: As media focuses on the election, Obama  implements most destructive plans behind the scenes.https://t.co/A"
TineCrane1|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
TineCrane1||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
SquishyBomb1|BushwackCA|-0.8109|0.295|0.705|0.0|"RT @BushwackCA: So if #Russia ""Hacked the US election"" then maybe #Hillary didn't win the popular vote. I would bet Russia would rather dea"
SFDoug|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
RobinSeaholm|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
rundiwala|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
rundiwala|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
DavidMoralee|youtube|-0.6908|0.289|0.711|0.0|"Arrogance &amp; Media Corruption, lost the DNC it's election, not #RussianInterference and still it continues.  https://t.co/wT30zOd14g"
foxmia1971|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
biggunz1965|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
keating_eleanor|LindaSuhler|-0.5574|0.247|0.753|0.0|RT @LindaSuhler: #FakeNews: CNN Shamed into Major Corrections on Ghana Election Storyhttps://t.co/czJezq4MlR
Get2KnowSaintJo|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
MarilynnePryor|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Huffaker3|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
pl8ofshrimp|jonhartmannjazz|0.0|0.0|1.0|0.0|@jonhartmannjazz @mmpadellan https://t.co/AtlfkHh7r1
pl8ofshrimp|petitions|0.0|0.0|1.0|0.0|@jonhartmannjazz @mmpadellan https://t.co/AtlfkHh7r1
LaCina52|Green_Footballs|-0.4767|0.124|0.876|0.0|"RT @Green_Footballs: Wondering what it would take for this country to say, ""Wait, this is wrong. We need to re-do this election."" Because h"
zeroinscw|cerenomri|0.0|0.0|1.0|0.0|"RT @cerenomri: Remember that one week during the election when the left was really, really concerned about anti-Semitism?They're supporti"
katgrneyes|CodeAud|0.0516|0.0|0.915|0.085|"RT @CodeAud: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous""https://t.co/NMnedgK9Fw"
katgrneyes|washingtonpost|0.0516|0.0|0.915|0.085|"RT @CodeAud: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous""https://t.co/NMnedgK9Fw"
strawberryheidi|mtracey|-0.25|0.095|0.905|0.0|"RT @mtracey: Dems' post-election lunacy closely resembles GOP birtherism, except in this case the paranoia is far more mainstream https://t"
strawberryheidi||-0.25|0.095|0.905|0.0|"RT @mtracey: Dems' post-election lunacy closely resembles GOP birtherism, except in this case the paranoia is far more mainstream https://t"
LaOkieKat|laurahollis61|-0.6486|0.238|0.762|0.0|"RT @laurahollis61: This whole ""Russians hacked the election"" story is the biggest load of crap since#Benghazi ""it-was-a-video."" Dems are d"
Iwillnotfall|POLITICOMag|0.0|0.0|1.0|0.0|"RT @POLITICOMag: For restive liberals, de Blasios re-election campaign will be a first big test in the Age of Trump: https://t.co/m3vww3bw"
Iwillnotfall|t|0.0|0.0|1.0|0.0|"RT @POLITICOMag: For restive liberals, de Blasios re-election campaign will be a first big test in the Age of Trump: https://t.co/m3vww3bw"
JamesDubhthaigh|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
jrountreeinc|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
Ah_muzings|SaintGimp|-0.659|0.197|0.803|0.0|RT @SaintGimp: The most frustrating thing about this Russia thing: there's no NEW info here. All the facts were known to the right people b
librarian5280|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
TaiRagan|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
MsScree|michaelianblack|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
MsScree|twitter|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
luanph0311|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
luanph0311|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
CragoDeb|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
nana5greatgrand|Irwin_Elaine|0.0|0.0|1.0|0.0|RT @Irwin_Elaine: @_0HOUR1 Here's a list of all the Foreign Governments who interfered in the last Pres election. I mean... donated to the
chulesee|LoisSmithers|-0.7096|0.222|0.708|0.071|RT @LoisSmithers: Read to end - NYT lets itself off the hook for its horrific coverage of election: Truth and Lies in the Age of Trump http
amansharmaaap|AamAdmiPartyFBD|0.5574|0.0|0.753|0.247|"RT @AamAdmiPartyFBD: On Municipality Election, #TeamFaridabad leadership @AbhashChandela &amp; @ranbirchandila clarifies that Party will not co"
CalypsoCats|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
JBarongen|citizentvkenya|-0.0516|0.14|0.671|0.189|RT @citizentvkenya: Gambias President Jammeh to challenge election loss at top court https://t.co/hKl09ZAe8B https://t.co/Xh77HXSiS1
JBarongen||-0.0516|0.14|0.671|0.189|RT @citizentvkenya: Gambias President Jammeh to challenge election loss at top court https://t.co/hKl09ZAe8B https://t.co/Xh77HXSiS1
leftcoastcoach|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
BonnieGranny|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
wvjoe911|JuddLegum|0.0|0.0|1.0|0.0|Trump adviser suggests election hacks were false flag operation by the Obama administration by @JuddLegum https://t.co/jVkA3eRwxB
wvjoe911|medium|0.0|0.0|1.0|0.0|Trump adviser suggests election hacks were false flag operation by the Obama administration by @JuddLegum https://t.co/jVkA3eRwxB
JeffCallahan75|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
GingerSpiceCin|ChicagoMGD|0.4767|0.0|0.853|0.147|RT @ChicagoMGD: @aliasvaughn @ezlusztig Reminder it isn't just the @CIA 16 other intelligence agencies had evidence of Russia's interferenc
Koustubh1|Being_Humor|-0.6249|0.186|0.814|0.0|RT @Being_Humor: So Shri @ArvindKejriwal ji made @SatyendarJain Satinder because Punjab election is coming. Worst kind of politics. Shamefu
Ostravaczech|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Ostravaczech||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
fbrown7628|neeratanden|0.0|0.0|1.0|0.0|@neeratanden @EricLiptonNYT @ScottShaneNYT @EricLichtblau @nytimes Get over it. Don't you offer more as a lib/dem?the election 4 1/2wks ago!
sguglie2|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
GamerOps|MaxAbrahms|-0.5106|0.136|0.864|0.0|RT @MaxAbrahms: The Twitter outrage over Russian interference in the election would be more credible if not spearheaded by Hillary fans loo
2crazy4books2|Sifill_LDF|0.0|0.0|1.0|0.0|@Sifill_LDF @ndylan1 https://t.co/UriwbWI930
2crazy4books2|petitions|0.0|0.0|1.0|0.0|@Sifill_LDF @ndylan1 https://t.co/UriwbWI930
snickerfritz04|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
e_revolutionist|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
melissa_sawyer|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
disgustedvoter2|Lee_in_Iowa|-0.5719|0.171|0.829|0.0|"RT @Lee_in_Iowa: Hey, @realDonaldTrump, in case you thought you actually ""won"" the election, no.Americans hate you. Oh well..... https://t"
disgustedvoter2||-0.5719|0.171|0.829|0.0|"RT @Lee_in_Iowa: Hey, @realDonaldTrump, in case you thought you actually ""won"" the election, no.Americans hate you. Oh well..... https://t"
clausen_ed|colinjones|0.3182|0.116|0.677|0.207|"RT @colinjones: You know, Im, like, a smart person. - Trump on criticism of his refusal of more regular intel briefings https://t.co/aGd"
clausen_ed|t|0.3182|0.116|0.677|0.207|"RT @colinjones: You know, Im, like, a smart person. - Trump on criticism of his refusal of more regular intel briefings https://t.co/aGd"
ALKCFA|stephenWalt|-0.4019|0.124|0.876|0.0|"RT @stephenWalt: Shocking that Russia tried to influence US election.  I mean, WE would NEVER interfere in another state's internal politic"
whaaf|scottwongDC|-0.34|0.112|0.888|0.0|"RT @scottwongDC: In rare bipartisan statement, McCAIN, GRAHAM, SCHUMER &amp; REED say reports of Russian interference in election ""should alarm"
phyzzycyst|Bill_Rhodes54|-0.3182|0.213|0.669|0.117|"RT @Bill_Rhodes54: #RussiaHacking is what you say when you:1) lose election2) realize ""popular vote"" means nothing3) Get humiliated by"
80sRetroPics|bbc|0.0|0.0|1.0|0.0|#Vintage #Retro #80s Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/BYThUsnLL8
SheilaSteger|HuffingtonPost|0.4939|0.083|0.728|0.189|RT @HuffingtonPost: These super PAC donors were able to hide their identities before the election https://t.co/J3NMv5ynDt https://t.co/Hyne
SheilaSteger|m|0.4939|0.083|0.728|0.189|RT @HuffingtonPost: These super PAC donors were able to hide their identities before the election https://t.co/J3NMv5ynDt https://t.co/Hyne
Smokyjo1|YouTube|0.0|0.0|1.0|0.0|CIA Splinter Group Calls For Overthrow Of Trump Election https://t.co/T488iiYWMG via @YouTube
Smokyjo1|youtube|0.0|0.0|1.0|0.0|CIA Splinter Group Calls For Overthrow Of Trump Election https://t.co/T488iiYWMG via @YouTube
DevilsGodson75|newcenturytimes|0.0|0.0|1.0|0.0|https://t.co/a94qZtoFZ5
PazyAmor53|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
InfoPasser|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
iTheHammer|JBurtonXP|0.6597|0.0|0.779|0.221|"RT @JBurtonXP: If Russia wanted to influence the election, they should've just donated millions to Hillary like all the respectable foreign"
kurt_cagle|twitter|0.4336|0.158|0.516|0.326|"Given the role the FBI played in the election, I share as hell trust the CIA more as an authority. https://t.co/MA8nzDjMD3"
SDReyley|ericgarland|0.0|0.0|1.0|0.0|RT @ericgarland: Do you tell America the day after the election that Russia spearfished all of our think tanks in brazen fashion?
ThomasKeown1|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
Pastapharian700|MtnMD|0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
Pastapharian700||0.0|0.0|1.0|0.0|RT @MtnMD: RT @asJBdorightthng: '94 SCOTUS:Mark v Stinson reversed state Sen election:2 officials knew R fraud-gv 2Dem opponent https://t.c
jamesmurphypdx|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
IslamophobiaLOL|barenakedislam|0.0|0.0|1.0|0.0|FLYING PIGS MOMENT from a far left writer at the New York Times: Election https://t.co/a2Xtae8A8r #islamophobia
BellaDawn01527|mabrams|0.0|0.0|1.0|0.0|"RT @mabrams: McCain, Graham, Schumer, Reed Joint Statement on Reports That Russia Interfered with the 2016 Election  https://t.co/sNuGY23cH1"
BellaDawn01527|armed-services|0.0|0.0|1.0|0.0|"RT @mabrams: McCain, Graham, Schumer, Reed Joint Statement on Reports That Russia Interfered with the 2016 Election  https://t.co/sNuGY23cH1"
GivingFace|youtube|-0.5423|0.32|0.552|0.127|The Truth About Fake News | Russia Hacked U.S. Election For Donald Trump? https://t.co/NJh3Gm6wjA
AsianAmeri4HRC|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
AsianAmeri4HRC|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
ChrisGaryL|LibertyTwoNews|-0.4767|0.171|0.829|0.0|RT @LibertyTwoNews: Sheryl Sandberg Says Fake News Did Not Sway Election | The Daily Caller https://t.co/GCIk9xhCDy  #breaking
ChrisGaryL|dailycaller|-0.4767|0.171|0.829|0.0|RT @LibertyTwoNews: Sheryl Sandberg Says Fake News Did Not Sway Election | The Daily Caller https://t.co/GCIk9xhCDy  #breaking
buffalogiu|igorvolsky|0.7845|0.0|0.711|0.289|RT @igorvolsky: Republicans used to love Congressional investigations. Will they support a probe into Russian hacking of the election? http
StateoftheInter|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
kountrykaye1257|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
JaneMoss08|jkarsh|0.4576|0.0|0.87|0.13|"RT @jkarsh: Given the CIA report about Russia influencing our election, this line from an @azcentral piece is very interesting. https://t.c"
JaneMoss08||0.4576|0.0|0.87|0.13|"RT @jkarsh: Given the CIA report about Russia influencing our election, this line from an @azcentral piece is very interesting. https://t.c"
marie_harl|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
marie_harl||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
bichonpawz|abc10|0.4404|0.101|0.671|0.228|'Make America Kind Again' signs in high demand even after election https://t.co/iwbAyeZdiC
PrincessBibiRF_|CarmineZozzora|0.0516|0.097|0.798|0.105|"RT @CarmineZozzora: Nothing like the CIA saving all their Russia ""secret assessment"" stuff up until after ""shoo-in"" Hillary lost the electi"
JRehling|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
PhyllisCopeland|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
boudreaulorrain|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
boudreaulorrain|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
SocialTweet509|_Makada_|-0.9081|0.383|0.617|0.0|RT @_Makada_: The same fake news media who said Iraq had weapons of mass destruction now claims Russia hacked our election. MSM are known l
fickles|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
fickles|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
cassroy|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
jodi_yoho|WeNeedTrump|-0.5413|0.155|0.845|0.0|RT @WeNeedTrump: Donald Trump's use of Twitter absolutely destroyed the mainstream media during this election. Will they ever learn? #MAGA
ginjasnappy|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
575haiku|adirado29|-0.5423|0.189|0.811|0.0|RT @adirado29: Moscow rules? CIA report raises troubling questions about Donald Trump's relationship with Russia https://t.co/wp0yNEhF4Q
575haiku|theage|-0.5423|0.189|0.811|0.0|RT @adirado29: Moscow rules? CIA report raises troubling questions about Donald Trump's relationship with Russia https://t.co/wp0yNEhF4Q
RebeccaSWH|scottwongDC|-0.34|0.112|0.888|0.0|"RT @scottwongDC: In rare bipartisan statement, McCAIN, GRAHAM, SCHUMER &amp; REED say reports of Russian interference in election ""should alarm"
PainePill|twitter|0.0|0.0|1.0|0.0|"These Yanks were open about foreign election intervention, unlike when the CIA has done it in Latin America. https://t.co/hVJ4F8WpFC"
virende19391800|cctvnews|-0.3612|0.161|0.839|0.0|RT @cctvnews: Donald Trump: CIA assessment of Russian interference in US election ridiculous https://t.co/faCCIwg7Ef
virende19391800|twitter|-0.3612|0.161|0.839|0.0|RT @cctvnews: Donald Trump: CIA assessment of Russian interference in US election ridiculous https://t.co/faCCIwg7Ef
charlescollier|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
lycoris_aurea|MrJamesonNeat|-0.6597|0.241|0.759|0.0|"RT @MrJamesonNeat: Read this comment, and sign the petition. In states where election fraud seems rampant lawsuits shoul... https://t.co/ms"
lycoris_aurea|twitter|-0.6597|0.241|0.759|0.0|"RT @MrJamesonNeat: Read this comment, and sign the petition. In states where election fraud seems rampant lawsuits shoul... https://t.co/ms"
Linda3717|jmsexton_|0.2263|0.079|0.794|0.127|"RT @jmsexton_: As Democrats demand probe over CIA election claim, GOP senators play politics. https://t.co/KNYgsIvWCx ~ @WashingtonPost htt"
Linda3717|washingtonpost|0.2263|0.079|0.794|0.127|"RT @jmsexton_: As Democrats demand probe over CIA election claim, GOP senators play politics. https://t.co/KNYgsIvWCx ~ @WashingtonPost htt"
mantalicious|ConsultDrSteve|0.0|0.0|1.0|0.0|"RT @ConsultDrSteve: BREAKING: Mitch McConnell Implicated In Russia/Trump Election Meddling, FBI Inquiry https://t.co/BVWtjsFLvW"
mantalicious|bipartisanreport|0.0|0.0|1.0|0.0|"RT @ConsultDrSteve: BREAKING: Mitch McConnell Implicated In Russia/Trump Election Meddling, FBI Inquiry https://t.co/BVWtjsFLvW"
therussophile|therussophile|0.0772|0.0|0.925|0.075|Secret Agenda: Are They Planning To Use Russian Interference As An Excuse To Invalidate Trumps ElectionVictory? https://t.co/pRjO9b7jPG
Top_Story_News|traffic|0.296|0.0|0.879|0.121|"Key GOP senators join call for bipartisan Russia election probe, even as their leaders remain mum https://t.co/KVgJjNSyWO"
mdurand1949|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
commentor2013|FBI|0.0|0.0|1.0|0.0|@FBI breaks with @CIA on Russia interference in U.S. election https://t.co/VlOlKLg6zE
commentor2013|thehill|0.0|0.0|1.0|0.0|@FBI breaks with @CIA on Russia interference in U.S. election https://t.co/VlOlKLg6zE
BenTurner15|nytimes|0.8442|0.0|0.637|0.363|"RT @nytimes: U.S. intelligence agencies have ""high confidence"" Russia acted covertly to help Trump in election, officials said https://t.co"
BenTurner15|t|0.8442|0.0|0.637|0.363|"RT @nytimes: U.S. intelligence agencies have ""high confidence"" Russia acted covertly to help Trump in election, officials said https://t.co"
SierranWolf|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
dimejibabalola|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
timothyworkman9|LindaSuhler|-0.2168|0.144|0.75|0.106|RT @LindaSuhler: Remember Obama's hot mic msg to Putin about flexibility after the election?What are they scared of? #RussianHackinghttps
d_a_keldsen|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
d_a_keldsen|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
NurseRatchets|DailyNewsBin|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
NurseRatchets|palmerreport|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
APendergast63|genebsperling|-0.5095|0.193|0.721|0.085|"RT @genebsperling: So at end of close election, FBI deeply hurt HRC based on no evidence, while CIA sat on clear evidence of Putin interfer"
jontalton|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
OurPowderDry|RBReich|-0.5719|0.179|0.821|0.0|@RBReich EC its Hillary.Thieves get stripped of ill-gotten goods  This cannot be turned over 2 Treasonous GOP. See  https://t.co/S2m37OCzm7
OurPowderDry|change|-0.5719|0.179|0.821|0.0|@RBReich EC its Hillary.Thieves get stripped of ill-gotten goods  This cannot be turned over 2 Treasonous GOP. See  https://t.co/S2m37OCzm7
ArdittoKime|PeterFosterALP|-0.4588|0.15|0.85|0.0|RT @PeterFosterALP: What a fizza.No wonder Australians are fed up with all the deceit of Malcolm Turnbulls fraudband https://t.co/ZEVqV
ArdittoKime|t|-0.4588|0.15|0.85|0.0|RT @PeterFosterALP: What a fizza.No wonder Australians are fed up with all the deceit of Malcolm Turnbulls fraudband https://t.co/ZEVqV
SimoneSmith3|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
_Carja|LampOlive|-0.8004|0.255|0.745|0.0|RT @LampOlive: We all knew Trump couldn't win without rigging the election. Getting Russia to do it is the worst Avenue to go.
sethmoulton|twitter|0.6808|0.0|0.797|0.203|"Proud to see so many #MA6 constituents ready to work for change. There is so much to do, and this election was a ca https://t.co/gHoHKmjkIO"
marclippincott|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
pankajtpatel|bleacherreport|0.0|0.0|1.0|0.0|"Doug Baldwin Comments on Donald Trump's Election, Inequality and More https://t.co/eOxC0XKA8b"
mau4682|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
HearMeRoar53881|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
CipollaKate|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
WhoFdTheStork|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
WhoFdTheStork||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
travel611|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
DestructiveChem|ReaganBattalion|0.1531|0.088|0.796|0.115|"RT @ReaganBattalion: Although liberals are hesitant to give him credit, Senator @MarcoRubio has been speaking about Russia meddling in our"
HerYin|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
HerYin||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
dmcobbphoto|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
mirakyz|ezlusztig|0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
mirakyz||0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
AziziOthmanMY|in|0.0|0.0|1.0|0.0|Trump says reports Russia helped him in U.S. election are 'ridiculous' https://t.co/KFWbV5URbY Trump says reports Russia helped him in U.S
hk_ravenclaw|PalmerReport|-0.4215|0.141|0.859|0.0|RT @PalmerReport: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day - https://t.co/TtRR8DcFBG
hk_ravenclaw|palmerreport|-0.4215|0.141|0.859|0.0|RT @PalmerReport: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day - https://t.co/TtRR8DcFBG
MiddletonSophia|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
JoshNoneYaBiz|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
azpat0|youtube|-0.7865|0.409|0.591|0.0|CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia https://t.co/UXIwN9I0nz
pakobserver|pakobserver|0.0|0.0|1.0|0.0|Romanian left seeks electioncomeback https://t.co/OH3uUCy2eu
BarboniMacaroni|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
BarboniMacaroni|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
caroljdavy|AdamsFlaFan|0.0|0.0|1.0|0.0|"RT @AdamsFlaFan: WAKE UP, AMERICA!!! Putin has interfered with our election and installed a puppet. We voted for Hillary. She leads trump b"
mike95465073|KellyannePolls|-0.7531|0.334|0.605|0.061|Conway calls CIA report on Russian election meddling laughable and ridiculous https://t.co/npA32dpk7k @KellyannePolls STUPID SKANK
mike95465073|washingtonpost|-0.7531|0.334|0.605|0.061|Conway calls CIA report on Russian election meddling laughable and ridiculous https://t.co/npA32dpk7k @KellyannePolls STUPID SKANK
trevordorn|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
mybodyGG|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
mybodyGG|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
poodbit499|twitter|-0.516|0.234|0.661|0.105|"Yes OBAMA hates BiBi so much he interfered w/Israels election &amp; tried to oust him,yet he's trying 2 BLAME Russia 4 https://t.co/nLCKRzIYaZ"
Saya_relativity|Khanoisseur|0.0|0.0|1.0|0.0|"RT @Khanoisseur: Looked at people in Whole Foods  line today and wondered ""how many of you thinking about the election rn?"" @michaelianblac"
Klayoven|Khanoisseur|-0.2263|0.087|0.913|0.0|RT @Khanoisseur: More new evidence that Comey tipped undecided voters toward Trump in last 2 weeks of the electionBiggest tamperer was th
againstabusesa|ewn|-0.3612|0.185|0.815|0.0|Trump says reports Russia helped him in US election are ridiculous https://t.co/tBfYF3JitO
crosa1988|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
sir_animesh_Ji|AmarUjalaNews|0.0|0.0|1.0|0.0|RT @AmarUjalaNews:  ''           https://t.co/7pU9fbxzk6#upelections
sir_animesh_Ji|amarujala|0.0|0.0|1.0|0.0|RT @AmarUjalaNews:  ''           https://t.co/7pU9fbxzk6#upelections
SnoopandWillie|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
SnoopandWillie|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
sallyodum|cnadnqt|0.1174|0.116|0.713|0.171|"RT @cnadnqt: @williesband @Greg_Palast @DrJillStein And, to be fair, if we don't fix these problems even a new election will be unfair and"
lesliern92|JeffCallahan75|0.25|0.105|0.752|0.143|@JeffCallahan75 how u figure? It's actually the KGB (Putin) that worries me. If Trump meant to be Pres. he can win a NEW election.
HelenEckard|Khanoisseur|0.5106|0.0|0.845|0.155|RT @Khanoisseur: .@LindseyGrahamSC Strong bipartisan statement on Russian meddling in election But you all need to also investigate FBI i
thinklightblue|nytopinion|0.0|0.0|1.0|0.0|RT @nytopinion: Why would President-elect Trump object to a thorough bipartisan probe into Russian meddling? https://t.co/zDopY4Hcs0 https:
thinklightblue|nytimes|0.0|0.0|1.0|0.0|RT @nytopinion: Why would President-elect Trump object to a thorough bipartisan probe into Russian meddling? https://t.co/zDopY4Hcs0 https:
sam_adjetey|NAkufoAddo|0.7269|0.0|0.775|0.225|"RT @NAkufoAddo: This morning, I attended the Ridge Church, Accra, with my family, to give thanks to the Lord for a peaceful election and gr"
MarkM447|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
MarkM447|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
carlastoneintl|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
pharmalady|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
lycoris_aurea|themattmcd|0.0|0.0|1.0|0.0|RT @themattmcd: Here is Mitch McConnell's office number:202-224-2541Call and ask why he kept us in the dark about foreign interference
AnneMcGibbs|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
BrianTDeegan|johnkennedyla|0.9098|0.0|0.511|0.489|Republican John Kennedy wins Louisiana senate race in runoff election https://t.co/y4EVIzEAiH - Congrats @johnkennedyla - great job!
BrianTDeegan|cnbc|0.9098|0.0|0.511|0.489|Republican John Kennedy wins Louisiana senate race in runoff election https://t.co/y4EVIzEAiH - Congrats @johnkennedyla - great job!
crosa1988|ElectoralCollge|-0.2846|0.203|0.702|0.095|@ElectoralCollge Russia rigged our election.Our true President is HRC.Dobt rob her.HRC can't b bought but Trump can https://t.co/lln2bjA22K
crosa1988|twitter|-0.2846|0.203|0.702|0.095|@ElectoralCollge Russia rigged our election.Our true President is HRC.Dobt rob her.HRC can't b bought but Trump can https://t.co/lln2bjA22K
JessMe757|technowizardry|0.0|0.0|1.0|0.0|RT @technowizardry: Did #Russia really hack the election?Please vote and RT!
ValkyrieHanna7|HardiesDazza|0.0|0.0|1.0|0.0|@HardiesDazza @JoyceSt14976939 @ANOMALY1 @KellyannePolls @realDonaldTrump https://t.co/G8tjpvsyYF
ValkyrieHanna7|newyorker|0.0|0.0|1.0|0.0|@HardiesDazza @JoyceSt14976939 @ANOMALY1 @KellyannePolls @realDonaldTrump https://t.co/G8tjpvsyYF
e_revolutionist|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
e_revolutionist|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
margie_sg|PrisonPlanet|-0.5106|0.191|0.809|0.0|"RT @PrisonPlanet: Post election riots: FAILED.Jill Stein recount: FAILED.Intimidation of EC members: FAILED.""Fake news"": FAILED.""Russia"
_mylesjames_|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
anesam98|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
anesam98|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
jjauthor|laurahollis61|-0.6486|0.238|0.762|0.0|"RT @laurahollis61: This whole ""Russians hacked the election"" story is the biggest load of crap since#Benghazi ""it-was-a-video."" Dems are d"
athada|youtube|0.582|0.169|0.522|0.309|"#PEOTUS admits #LockHerUp was gimmick: ""Forget it. That plays great before the election. Now, we dont care, right?"" https://t.co/bgaendjktD"
AldoKaz|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
AldoKaz|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
eddie736|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
eddie736|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
wrdybrd|jameshamblin|0.0|0.0|1.0|0.0|RT @jameshamblin: So people believe a pizza place is a government sex ring but fancy themselves too savvy to look into Russian election int
azpat0|YouTube|0.6124|0.0|0.688|0.313|I liked a @YouTube video https://t.co/u0TS48IRxY Maximum Alert: Rogue CIA Working to Overthrow Trump Election
azpat0|youtube|0.6124|0.0|0.688|0.313|I liked a @YouTube video https://t.co/u0TS48IRxY Maximum Alert: Rogue CIA Working to Overthrow Trump Election
riverqueen|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
daquick07|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
hotmerthanyou|swin24|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
hotmerthanyou|thedailybeast|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
Dinosgurl|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: Also, there must be investigation of Comey @FBI. That he could know this &amp; decide to break all history to interfere w/"
sbca80|amjoyshow|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
sbca80|t|0.7291|0.0|0.746|0.254|RT @amjoyshow: .@MCFAUL tells #AMJoy it's looking very clear that #Russia has meddled with our election. RETWEET TO AGREE https://t.co/n3RH
CatherineLucer4|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Backstorymom1|linkis|-0.4215|0.286|0.714|0.0|Worries deepen about Russia's involvement in election https://t.co/iTKvOLuZr6
LisainPA|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
cturtle31|LindseyThiry|0.3612|0.0|0.762|0.238|.@LindseyThiry Looks like a @HillaryClinton rally right before the election.
RiskyLiberal|bryanbehar|0.0772|0.18|0.631|0.189|RT @bryanbehar: We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure justice
ginalove3232|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
bettyonline011|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
veve4heart|politicususa|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
veve4heart|twitter|0.4019|0.0|0.876|0.124|RT @politicususa: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co/m
primosbaby|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
RGBennettJr89|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
MaelinnHughes|leahmcelrath|0.7088|0.081|0.623|0.296|@leahmcelrath Same here. We must do everything we can to stop. Please sign petition at https://t.co/HcqLIIb4WN Hoping it will help! RTplease
MaelinnHughes|petitions|0.7088|0.081|0.623|0.296|@leahmcelrath Same here. We must do everything we can to stop. Please sign petition at https://t.co/HcqLIIb4WN Hoping it will help! RTplease
rugratfarm|abctweet100|0.0|0.0|1.0|0.0|RT @abctweet100: Let It Sink In-The Evidence is OVERWHELMING that Russia Interfered With Our Election #ElectoralCollege #MoralElectors #fai
jess_sandhu|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
imanewman442|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
GermanoDottori|latimes|-0.0258|0.144|0.719|0.138|RT @latimes: Prominent senators say Russian election interference should alarm all Americans https://t.co/5QprDsvyoi https://t.co/SuFzJ25R0b
GermanoDottori|latimes|-0.0258|0.144|0.719|0.138|RT @latimes: Prominent senators say Russian election interference should alarm all Americans https://t.co/5QprDsvyoi https://t.co/SuFzJ25R0b
cjstrickling|Moo57556470|-0.4943|0.2|0.714|0.086|"RT @Moo57556470: If Americans cannot trust its Congress, its FBI &amp; certainly its PEOTUS, how can we repair the damages absent A NEW ELECTIO"
randypitler|nsroundtable|-0.4019|0.119|0.881|0.0|@nsroundtable @ann_nooner @davidfrum @AlecMacGillis It is based on how this election went. What proof do you have that it was hacked?
dg2wright|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
trex9123|NPR|-0.7003|0.234|0.766|0.0|"@NPR @jasunmark I say this as $ a day member,but NPR's coverage of election this year just as bad as CNN's.Complete lack of proportionality."
LikusPJ|starfirst|-0.2003|0.107|0.893|0.0|RT @starfirst: Demand An Audit Of The 2016 Presidential Election - Sign the Petition! https://t.co/VPAVYiDzlX via @Change
LikusPJ|change|-0.2003|0.107|0.893|0.0|RT @starfirst: Demand An Audit Of The 2016 Presidential Election - Sign the Petition! https://t.co/VPAVYiDzlX via @Change
JessesLaw|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
JessesLaw||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
johnnyt74|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
LitLat|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
msjbe20a|buffaloon|0.2732|0.0|0.861|0.139|RT @buffaloon: Russia's Interference in This Election Should Not Be a Surprise https://t.co/HhshcPRbC4 via @Esquire
msjbe20a|esquire|0.2732|0.0|0.861|0.139|RT @buffaloon: Russia's Interference in This Election Should Not Be a Surprise https://t.co/HhshcPRbC4 via @Esquire
smegmalomaniac|cliffordlevy|0.0|0.0|1.0|0.0|"RT @cliffordlevy: The facts: since the election, @nytimes has seen a surge in new digital subscriptions, 6 times our normal pace https://t."
smegmalomaniac||0.0|0.0|1.0|0.0|"RT @cliffordlevy: The facts: since the election, @nytimes has seen a surge in new digital subscriptions, 6 times our normal pace https://t."
__solodolo__|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
__solodolo__||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
MrsBodie2|rwindrem|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
MrsBodie2|nbcnews|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
maewest80|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
DssdentAggrssor|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
TNChick67|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
TNChick67|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
hangthebankers|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
JamesAThomas67|latimes|0.2023|0.0|0.878|0.122|Trump faces first significant post-election pushback from Republicans over CIA report on Russia https://t.co/vhKmkJdUrU
BonnieGranny|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
annabelslil|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
joe_nca|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
PetsVoteToo|LauraBenanti|0.6669|0.143|0.604|0.253|RT @LauraBenanti: Don't let Trumps twitter rants distract from the real news: THE RUSSIANS INTERVENED IN OUR ELECTION TO HELP TRUMP WIN. #r
jkumac|PolitiFact|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
jkumac|t|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
Xaniatube|xaniatube|-0.1531|0.118|0.882|0.0|"New video: Morning Joe Host: Hillary Censored Us, Interfered In Election - https://t.co/B9SqLksyFU #XaniaTube"
PaceSociety|MyHarmReduction|0.0|0.0|1.0|0.0|RT @MyHarmReduction: A NYTimes article of Self-Care- buzzword or real therapeutic tool? https://t.co/8dFVQNZoRb
PaceSociety|nytimes|0.0|0.0|1.0|0.0|RT @MyHarmReduction: A NYTimes article of Self-Care- buzzword or real therapeutic tool? https://t.co/8dFVQNZoRb
snobbygirl17|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
PSW101|StrangeLondon|-0.7351|0.341|0.659|0.0|RT @StrangeLondon: The Gambia: troops deployed to streets as president rejects election defeat https://t.co/E8pR35WmOb
PSW101|theguardian|-0.7351|0.341|0.659|0.0|RT @StrangeLondon: The Gambia: troops deployed to streets as president rejects election defeat https://t.co/E8pR35WmOb
SoNortori_us|Complex|0.0516|0.192|0.604|0.203|"@Complex 1st Trump wins the election, now Dom Torito betrays his family #ThankForNothing2016"
dbergg|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
nuggiano1|Miami4Trump|0.368|0.129|0.684|0.187|RT @Miami4Trump: Hillary Is FILLED WITH GLEE Because WaPo Is Pushing Her Delusional Conspiracy Theory About Russia Hacking Our Election  #
TheOralBuffet|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
DavidWa39715864|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Geniusbastard|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
atomicrocketpop|FTI_US|0.6705|0.0|0.744|0.256|RT @FTI_US: #Zahn: We think Trumps election could provide a slight boost to the United Kingdoms #Brexit negotiations. https://t.co/NT6mE5
atomicrocketpop|t|0.6705|0.0|0.744|0.256|RT @FTI_US: #Zahn: We think Trumps election could provide a slight boost to the United Kingdoms #Brexit negotiations. https://t.co/NT6mE5
SOUTHERNjamespb|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
PegDelp|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
PegDelp|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
thenotsohotmess|guardiannews|0.0|0.0|1.0|0.0|RT @guardiannews: Romania's left takes big lead in parliamentary election - exit polls https://t.co/UTA3SGdL1N
thenotsohotmess|theguardian|0.0|0.0|1.0|0.0|RT @guardiannews: Romania's left takes big lead in parliamentary election - exit polls https://t.co/UTA3SGdL1N
TomMBell1|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
dgdocter12|60Minutes|0.2718|0.093|0.772|0.135|RT @60Minutes: .@netanyahu says Israel has never been in a better place; part of his optimism relates to the election of Trump https://t.co
dgdocter12|t|0.2718|0.093|0.772|0.135|RT @60Minutes: .@netanyahu says Israel has never been in a better place; part of his optimism relates to the election of Trump https://t.co
thewrightkansan|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
thewrightkansan||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
benonebo|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
benonebo|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
NakedSmBiz|hwcdn|0.296|0.0|0.833|0.167|Five small business experts share their post-election observations and recommendations https://t.co/QDctL5l18S https://t.co/cdZI5NmMcN
LikusPJ|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
zitab|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
JB_Hilterman|sea329|-0.7964|0.384|0.616|0.0|"RT @sea329: @DRUDGE_REPORT Hillary cheated, rigged the election and spent all that money and still lost "
whaaf|greenhousenyt|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
whaaf|t|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
clintonfein|JustinRaimondo|-0.4497|0.134|0.866|0.0|"@JustinRaimondo For a sec I thought you meant investigate renegade FBI agents involved in election tampering, but forgot you'd lost the plot"
TheWhiteNite83|TheFlightMike|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
TheWhiteNite83|twitter|0.0|0.0|1.0|0.0|RT @TheFlightMike: BREAKING: Tim Tebow and Johnny Manziel to run against Donald Trump in 2020 Presidential Election. https://t.co/eK499g6UD7
cussetabraswell|wonderfullone|0.0|0.0|1.0|0.0|RT @wonderfullone: Trump: It's 'Ridiculous' To Think Russia Intervened In The Election On My Behalf https://t.co/aQXguJxNsR
cussetabraswell|linkis|0.0|0.0|1.0|0.0|RT @wonderfullone: Trump: It's 'Ridiculous' To Think Russia Intervened In The Election On My Behalf https://t.co/aQXguJxNsR
curtoUSMC|BreitbartNews|-0.8959|0.34|0.66|0.0|"@BreitbartNews So bad, there has to be others turning this unfunny CRAP off besides me! My choice are videos of celebs crying over Election!"
Isabellarowling|ezlusztig|0.296|0.089|0.732|0.179|"@ezlusztig @Coreybez1 Well, since nothing was done to stop Trump before election, at least let the truth take Trump down after."
livetweettweet|MrJamesonNeat|-0.6597|0.231|0.769|0.0|RT @MrJamesonNeat: In states where election fraud seems rampant lawsuits should be filed to disqualify Trump electors @tribelaw @lessig htt
PoliticalBee|aliasvaughn|-0.3597|0.102|0.898|0.0|"RT @aliasvaughn: 9. So stop trying with ""oh they just ""tried to influence"" the election"" and start realizing that what we're dealing with i"
rickhasen|electionlawblog|-0.0772|0.091|0.909|0.0|#ELB; Sorry But Alleged Russian Influence in Presidential Election Wont Lead to a Do-Over https://t.co/qRyNjiCXmh
mirakyz|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/4TnN8g6MGt https://t."
mirakyz||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/4TnN8g6MGt https://t."
rphawg3150|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
DoloresWells20|20committee|0.7269|0.0|0.775|0.225|RT @20committee: Honest investigation of what Putin &amp; his spies did with our election this year will reveal truths that are deeply uncomfy
tom_luu|thehill|0.0|0.0|1.0|0.0|@thehill 2016 Election Recap: https://t.co/bLhh9FmlTl
tom_luu|twitter|0.0|0.0|1.0|0.0|@thehill 2016 Election Recap: https://t.co/bLhh9FmlTl
msjbe20a|buffaloon|-0.0516|0.162|0.684|0.154|"RT @buffaloon: Supreme Court: Election Can Be Invalidated Due To Massive Fraud, Install Opponent (DETAILS) https://t.co/eVFRhQtFgM via @Bip"
msjbe20a|bipartisanreport|-0.0516|0.162|0.684|0.154|"RT @buffaloon: Supreme Court: Election Can Be Invalidated Due To Massive Fraud, Install Opponent (DETAILS) https://t.co/eVFRhQtFgM via @Bip"
FrankNatale2|DrJillStein|0.0|0.0|1.0|0.0|"RT @DrJillStein: We expect bank tellers to double-check money before handing it to us. Let's double-check election results, too. #Recount20"
LalaFox4|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Gradebooks|PrankInvasion|0.5719|0.0|0.764|0.236|RT @PrankInvasion: Who else is happy this election is almost over? #voted #ElectionDay
2ALAW|LeahR77|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
2ALAW|t|0.0772|0.0|0.942|0.058|RT @LeahR77: Democrats Graham &amp; McCain Will Head Probe Into So Called Russian Influence Of Election &gt; Seems They Want WW3 https://t.co/JNhj
JonRuhe|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
AscanioMatt|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
AscanioMatt|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
lovemrpibb2|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/mEIzELKuVz https://t."
lovemrpibb2||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/mEIzELKuVz https://t."
aelmenhurst|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
logicalwing|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
logicalwing|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
MntsofWv|tteegar|-0.5242|0.232|0.67|0.098|RT @tteegar: BREAKING #RussianHackers made Hillary screech like an old crabby grandma &amp; lose the election!Nobody should be fooled! #Fak
daquick07|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
I_am_Mutated|Slate|-0.6544|0.172|0.828|0.0|"@Slate Election meddling? Oh you mean those leaks that proved DNC was the ones ""hacking"" &amp; stealing election by controlling media? Darn!..."
UnlikelyLass|twitter|0.8885|0.0|0.588|0.412|"They won the election, Rich. They got theirs, why would they care about the rest of us? https://t.co/VXlpKDQvI3"
librab103|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
petatusa|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Chaparro916|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
DocHoliday89|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
C2017DebouCracy|twitter|-0.2732|0.189|0.811|0.0|"#PrimaireDroite:https://t.co/89lIZUilj2 The election was stolen, but not by... https://t.co/F9XNsZGSCr https://t.co/yWHEDz2wP9"
RobbieLoucks|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
aintlifegrand99|jillybeans1203|-0.2144|0.112|0.811|0.077|RT @jillybeans1203: I should be surprised it took this crazy election for people to realize you shouldn't believe everything you read on th
mmdornconsult|thehill|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
mmdornconsult|twitter|-0.4201|0.202|0.798|0.0|"RT @thehill: Biden: Trump ran ""most vicious"" campaign I've ever seenhttps://t.co/60eCL3owHK https://t.co/rRCW6OVCmR"
takinyera|ericgarland|0.0|0.0|1.0|0.0|RT @ericgarland: Do you tell America the day after the election that Russia spearfished all of our think tanks in brazen fashion?
bchek833|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
Tracy_Mack|CaptainsLog2016|-0.4019|0.144|0.856|0.0|"RT @CaptainsLog2016: After election results are reversedTrumpkins will scream civil warThat's coolWe'll have Gov, police, &amp; American"
passionlaw|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
passionlaw|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
lipchikphoto|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
EmilyWA98498|thehill|-0.34|0.13|0.87|0.0|"RT @thehill: Bipartisan group of senators say Russian interference in the election should ""alarm every American""https://t.co/rypjh7XDrf ht"
EmilyWA98498|thehill|-0.34|0.13|0.87|0.0|"RT @thehill: Bipartisan group of senators say Russian interference in the election should ""alarm every American""https://t.co/rypjh7XDrf ht"
1984infoseeker|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
B_L_Mencken|twitter|-0.3472|0.125|0.808|0.067|"#Treason You can't  forget #JamesComey &amp; the shame he brought on himself, the FBI &amp; the nation. He emerges from the https://t.co/uAWdu8BeK9"
coleyhiles1|Melodic_prog|-0.5267|0.274|0.598|0.128|"Eh hem, who cares if a foreign nation hacked our election? You must hate this country @Melodic_prog @vicenews"
takief|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
doula_theou|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
dynamex|thehill|0.0|0.0|1.0|0.0|FBI breaks with CIA on Russia interference in U.S. election https://t.co/Gk6WQTFO1u
cattsmall|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
quest23blue|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
CerulloElaine|WeNeedTrump|-0.4522|0.129|0.871|0.0|"RT @WeNeedTrump: So the left cries about Russia allegedly interfering with our election. Yet, millions were donated to the Clinton Foundati"
LRD90|JuddLegum|0.0|0.0|1.0|0.0|RT @JuddLegum: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/oRUPSkz7NV https:
LRD90|medium|0.0|0.0|1.0|0.0|RT @JuddLegum: Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/oRUPSkz7NV https:
croesus2009|newsbusters|0.0|0.0|1.0|0.0|CNN's Robert Baer: We Should Have Another Election https://t.co/IpUos82miy
odinsbeer|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
GHFiii|PGEddington|-0.3642|0.277|0.564|0.159|RT @PGEddington: Americas most notorious intelligence agency says #Election2016 was hacked. The proper response: https://t.co/ASpIV1rpfn
GHFiii|medium|-0.3642|0.277|0.564|0.159|RT @PGEddington: Americas most notorious intelligence agency says #Election2016 was hacked. The proper response: https://t.co/ASpIV1rpfn
KoRickZenz|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
LALakerSh0rty|Opa001|-0.4588|0.2|0.8|0.0|RT @Opa001: Gambia leader Yahya Jammeh to contest election defeat in court https://t.co/8VFTy07KKE
LALakerSh0rty|bbc|-0.4588|0.2|0.8|0.0|RT @Opa001: Gambia leader Yahya Jammeh to contest election defeat in court https://t.co/8VFTy07KKE
Stevenb2|MissLizzyNJ|-0.952|0.53|0.47|0.0|"RT @MissLizzyNJ: #ImStillNotOver the fact that I lost the election because I'm a lying criminal and America hates me, so I'll blame fake ne"
amorganfloyd13|armed-services|0.0|0.0|1.0|0.0|https://t.co/hfS9810Aj4 https://t.co/UyJSMkRlJk
RedApplePol|npr|0.0|0.0|1.0|0.0|President Obama Orders 'Full Review' Of Hacking During 2016 Election : #TrumpRussia#notmypresident #CNNGetItRight  https://t.co/g8rXfMzfVz
ZoranTaylor|sarahclazarus|0.3182|0.0|0.901|0.099|RT @sarahclazarus: We'll know for sure the Russians were involved if we look into the election and find a smaller election right inside
WoodlandsTrudy|Stevenwhirsch99|0.5659|0.0|0.811|0.189|RT @Stevenwhirsch99: About a month and a half ago Obama told America elections couldn't be hacked. Now he's saying our election has been ha
yugvaniworld|in|0.0|0.0|1.0|0.0|Trump says reports Russia helped him in U.S. election are 'ridiculous' https://t.co/ktmoTqCyNI
wendellshaw5|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
Ava386|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ProfCAnderson|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
Kmich718|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
Kmich718|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
Deejdelo|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
dg2wright|LeahR77|0.1531|0.11|0.758|0.133|RT @LeahR77: Lets Talk Foreign Govts Influencing An Election &amp; Bonus Getting Uranium &amp; Weapons Deals From SOS HRC For #FakeNews #Russians
vquagliana|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
NrIsodera|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
NelsonForTruth|PeacefulChrist|0.0|0.0|1.0|0.0|RT @PeacefulChrist: @realDonaldTrump @ReiserWilliam @michaelmeans49 @MiceeMouse @perossmeisl #Election #election2016 recount 80 #Polling ma
Lolly_Jean|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
Sisterwriter|washingtonpost|0.296|0.0|0.879|0.121|"Key GOP senators join call for bipartisan Russia election probe, even as their leaders remain mum https://t.co/Hf7fqXR27u"
rcdubose|igorvolsky|0.7695|0.049|0.717|0.234|"RT @igorvolsky: The GOP position on foreign countries trying to rig our election seems to be: WE'RE OKAY WITH IT, AS LONG AS WE WIN."
cat_1012000|MaydnUSA|-0.4019|0.119|0.881|0.0|"RT @MaydnUSA: When Sony was hacked, the FBI immediately produced evidence. Anyone seen any actual evidence of election hack by Russia?Did"
HeyNikki1|jalloyd4|0.7579|0.0|0.683|0.317|"RT @jalloyd4: #CIA concludes Russia interfered to help Trump win #election, say reports @guardian https://t.co/Fj70RFINl4 #TheResistance"
HeyNikki1|theguardian|0.7579|0.0|0.683|0.317|"RT @jalloyd4: #CIA concludes Russia interfered to help Trump win #election, say reports @guardian https://t.co/Fj70RFINl4 #TheResistance"
cikoontz|PolitiFact|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
cikoontz|t|-0.296|0.121|0.879|0.0|RT @PolitiFact: False: Priebus falsely claims no conclusive report whether Russia tried to influence election. @MeetThePress https://t.co/Y
ChrisRiley001|cnn|0.0|0.0|1.0|0.0|We need an investigation into Russian interference in our election. https://t.co/SStk9kUudb
ggindc|scarylawyerguy|0.2052|0.08|0.805|0.114|"RT @scarylawyerguy: Special Benghazi Cmte after 7 other invests turned up nothing is ok, finding out if Russia interfered w/our election is"
tom_luu|PJStrikeForce|0.0|0.0|1.0|0.0|@PJStrikeForce 2016 Election Recap: https://t.co/bLhh9FmlTl
tom_luu|twitter|0.0|0.0|1.0|0.0|@PJStrikeForce 2016 Election Recap: https://t.co/bLhh9FmlTl
odom_1|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
erichstrat|howiewolf|0.0772|0.0|0.933|0.067|RT @howiewolf: Number of Congressional hearings on Benghazi: 33.Number of Congressional hearings on Russian efforts to influence our elec
Tuffelhund2003|Meow1113|0.0|0.0|1.0|0.0|"@Meow1113 @washingtonpost He'll get 4 years o correct BHO last 8, then we do another election."
cball47|FoxNewsSunday|0.0|0.0|1.0|0.0|RT @FoxNewsSunday: Coming up on #FNS -- @realDonaldTrump describes what went through his mind on election night. https://t.co/tJ7myY6Sxk
cball47|twitter|0.0|0.0|1.0|0.0|RT @FoxNewsSunday: Coming up on #FNS -- @realDonaldTrump describes what went through his mind on election night. https://t.co/tJ7myY6Sxk
ralphbod|igorvolsky|0.7845|0.0|0.711|0.289|RT @igorvolsky: Republicans used to love Congressional investigations. Will they support a probe into Russian hacking of the election? http
withrainyeyes|justbraden|-0.4404|0.172|0.828|0.0|RT @justbraden: Biggest tragedies of 2016:1. Harambe (RIP)2. Presidential Election3. Me not getting a text back
mattiOgreen|leahmcelrath|-0.3412|0.112|0.888|0.0|RT @leahmcelrath: NYTimes Editorial Board takes a stand &amp; even calls Trump out for not supporting an investigation into Russia hackinghttp
maryverobeach|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Michaelleschmid|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
Michaelleschmid|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
takinyera|ericgarland|-0.296|0.099|0.901|0.0|RT @ericgarland: Do you come out the day after this totally weird-smelling abomination of an election with all its technical difficulties?
LauraK205|LOLGOP|0.25|0.058|0.846|0.096|RT @LOLGOP: This election is like if A Christmas Carol ended with Scrooge getting a giant tax break paid for by cutting Tiny Tim off Medica
JackRoss061485|ScottMcConnell9|-0.5994|0.157|0.843|0.0|"RT @ScottMcConnell9: Election comes down to victory for: open borders, showdown w. Russia, ""free"" trade, war on cops or victory for bombast"
HarishC60347066|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
valeyrie47|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/mEIzELKuVz https://t."
valeyrie47||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/mEIzELKuVz https://t."
travel611|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
Daneuntamed|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
RobinWood|thehighsign|-0.1027|0.065|0.935|0.0|RT @thehighsign: If only someone had tried to warn us about this Russian hacking business _before_the election. At a podium. During a debat
Jjcruz2|twitter|0.0|0.0|1.0|0.0|Ediwow! Kayo na ung malinis na naulol nun election...  https://t.co/ZQ29EAQ3g3
Naijai3|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
TheKStainback|ezlusztig|0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
TheKStainback||0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
ayawill|ChrisCuomo|0.4767|0.0|0.83|0.17|RT @ChrisCuomo: Trump team still defending win. start defending US cyber security. Election over. Putin should be target but he isn't. Why?
Charonronn|joanneprada|-0.5719|0.381|0.619|0.0|RT @joanneprada: 2016 election: the ultimate scam
triniellis|mcw0530|-0.0108|0.112|0.778|0.11|@mcw0530 @mikd33 @ckkoch3 @JhoniiAlmeida note I didn't lose anything. America lost the election as Russia with Wikileaks hijacked it.
mccuebillie|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
mccuebillie||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
GS__User|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
marcylauren|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
Supertoaste|ECrowleyBooks|-0.6808|0.301|0.699|0.0|"RT @ECrowleyBooks: @politico He attacks everyone, except the foreign power that hacked our election. https://t.co/j0eDBlrYgD"
Supertoaste|twitter|-0.6808|0.301|0.699|0.0|"RT @ECrowleyBooks: @politico He attacks everyone, except the foreign power that hacked our election. https://t.co/j0eDBlrYgD"
grhodes123|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
grhodes123|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
777Francejacque|V_of_Europe|0.1027|0.162|0.614|0.224|RT @V_of_Europe: Italian Eurosceptics furious over MPs trying to secure pension boost in General Election https://t.co/8ppYHixKwN https://
777Francejacque|express|0.1027|0.162|0.614|0.224|RT @V_of_Europe: Italian Eurosceptics furious over MPs trying to secure pension boost in General Election https://t.co/8ppYHixKwN https://
NelsonForTruth|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
lycoris_aurea|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
lycoris_aurea||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
xocolleenxoxo|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
johnnyt74|michaelianblack|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
johnnyt74|twitter|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
melvyl|PastVox|0.7839|0.0|0.744|0.256|"RT @PastVox: 1968: Election analysis from Vox's Tate Silver ""Dem hopeful Robert Kennedy would've beat Nixon by 3 points were he not killed"
DeelightRI|MystryGAB|0.6124|0.0|0.762|0.238|RT @MystryGAB: @SenatorIsakson Please support the investigation into Russia's involvement in election. This is not partisan. Americans need
SOFTNOCTIS|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
SOFTNOCTIS|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
life_benefit|BrittPettibone|-0.4588|0.13|0.87|0.0|"RT @BrittPettibone: #ImStillNotOver the fact that, after being savaged by WikiLeaks during the U.S. Election, the MSM still believes it has"
icenite|DannyZuker|0.7184|0.0|0.76|0.24|"RT @DannyZuker: PATRIOT TEST:  If you're cool with Russia meddling with our election because your candidate won, you're not a patriot. Also"
whatistheimpact|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Dylan_Sandas|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
Dylan_Sandas|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
fixedopsjack|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
fixedopsjack|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
LoriRLopez|nytimes|-0.4767|0.171|0.829|0.0|Major #denial Trump Links C.I.A. Reports on Russia to Democrats Shame Over Election https://t.co/Ox5mtwPwv5 #NotMyPresident #StillWithHer
Donna_DHKBB|scoootchover|0.0|0.0|1.0|0.0|RT @scoootchover: @JoyAnnReid They have my vote to re-vote. #LetTheTruthWin #StillWithHerhttps://t.co/laBzxzoyUR
iTheHammer|JBurtonXP|-0.4019|0.124|0.876|0.0|"RT @JBurtonXP: Always remember that by ""hacked the election,"" these people mean ""released 100% authentic documents that showed real Democra"
ce06799|tgreene319|0.0|0.0|1.0|0.0|RT @tgreene319: Let's review. CIA says Russian hackers interfered w election. Russia says they didn't. Trump doesn't believe CIA &amp; instead
Collette_AZ|mtracey|-0.3595|0.098|0.902|0.0|@mtracey No to a new election w/out all 50 states voter id laws. W/NOT take hrs again out of workday &amp; spend Billions . Elections OVER!
Bannreyes|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
StevenNantz|PattyMurray|0.6124|0.0|0.75|0.25|"@PattyMurray Yes. Senator, please insist on a bipartisan investigation of Russian intervention in the 2016 U.S. presidential election."
postofficetruth|csmonitor|0.2023|0.0|0.886|0.114|RT @csmonitor: Obama's top counterterrorism adviser Lisa Monaco says key stakeholders need fuller answers. https://t.co/qXbRUYNHcQ
postofficetruth|csmonitor|0.2023|0.0|0.886|0.114|RT @csmonitor: Obama's top counterterrorism adviser Lisa Monaco says key stakeholders need fuller answers. https://t.co/qXbRUYNHcQ
kturet|SamWangPhD?|-0.4215|0.259|0.741|0.0|"The election just broke you, didn't it @SamWangPhD? https://t.co/f9zqmzIE9Q"
kturet|twitter|-0.4215|0.259|0.741|0.0|"The election just broke you, didn't it @SamWangPhD? https://t.co/f9zqmzIE9Q"
contrarian_prag|ejenk|0.7906|0.0|0.696|0.304|RT @ejenk: I saw a video of Russians cheering on the rooftops in New Jersey when Trump won the election.
SimplementeSole|2crazy4books2|0.0|0.0|1.0|0.0|RT @2crazy4books2: @Serpentine202 The CIA has proof. GOP conspired to suppress. https://t.co/UriwbWI930
SimplementeSole|petitions|0.0|0.0|1.0|0.0|RT @2crazy4books2: @Serpentine202 The CIA has proof. GOP conspired to suppress. https://t.co/UriwbWI930
OutHouseAtty|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
OutHouseAtty|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
Sailfish157|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
Sailfish157|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
tahino1|penultimatepen|0.4019|0.0|0.876|0.124|RT @penultimatepen: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co
tahino1|t|0.4019|0.0|0.876|0.124|RT @penultimatepen: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co
Sheptacular|igorvolsky|-0.4019|0.13|0.87|0.0|RT @igorvolsky: GOP Congressmembers react to news that Russia hacked election to aid Trump 1 called for investigations1 dismissed it301
longgoneblond|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
longgoneblond||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
StoneColdChik|rt|-0.4939|0.176|0.824|0.0|this is hillary obama mccain graham burr and this administration attempting to steal the election https://t.co/FsC7FQ1FEG
ChrisZametz|1Kimsey|0.2057|0.0|0.878|0.122|RT @1Kimsey: Why not? Jeh Johnson didn't hesitate to hack during GA election. https://t.co/vri97ni1yR
ChrisZametz|twitter|0.2057|0.0|0.878|0.122|RT @1Kimsey: Why not? Jeh Johnson didn't hesitate to hack during GA election. https://t.co/vri97ni1yR
angielashaye|TheRevAl|0.6416|0.057|0.762|0.181|@TheRevAl March on Washington? Really? 2 mths post election?Think it's time Black America gets some tough love. Tell us to take our medicine
ButtaSW|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
reasonandlogic|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
DamianSalizar|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
DamianSalizar|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
MartyTruthHurts|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
MartyTruthHurts||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
JeramySinopoli|YouTube|0.0|0.0|1.0|0.0|Ex-CIA operative calls for new election https://t.co/x2PkDaHikd via @YouTube
JeramySinopoli|youtube|0.0|0.0|1.0|0.0|Ex-CIA operative calls for new election https://t.co/x2PkDaHikd via @YouTube
cikoontz|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
cikoontz|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
Katie_Toledo1|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
jrountreeinc|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
kencf0618|SilverbearHeart|0.2682|0.0|0.901|0.099|RT @SilverbearHeart: After Trump's election ...... Russian influence in the GOP is systemic and more far reaching than Trump https://t.co/t
kencf0618|twitter|0.2682|0.0|0.901|0.099|RT @SilverbearHeart: After Trump's election ...... Russian influence in the GOP is systemic and more far reaching than Trump https://t.co/t
zoomie2012|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
LoriLevin|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
Yombe|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
leoluminary|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
leoluminary|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
MarieMurcelle1|conlimonisal|0.0|0.0|1.0|0.0|"RT @conlimonisal: @Greg_Palast I don't understand why Hillary hasn't requested recount,considering all of the election tampering allegation"
naretevduorp|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ZTOESQ|cushbomb|0.128|0.126|0.69|0.184|RT @cushbomb: If a failing petrooligrachy like Russia can determine the outcome of a presidential election it's fair to say America is not
HigginsSusan2|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
aandrewsaz|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
davisindy|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
postofficetruth|blckdetroit|0.0772|0.108|0.769|0.123|"RT @blckdetroit: Obama Administration Orders Probe Into Russia Election Hack Charges: Lisa Monaco, Homeland Security and https://t.co/msxs"
postofficetruth|t|0.0772|0.108|0.769|0.123|"RT @blckdetroit: Obama Administration Orders Probe Into Russia Election Hack Charges: Lisa Monaco, Homeland Security and https://t.co/msxs"
DiscoPotential|michaelianblack|0.0|0.0|1.0|0.0|"@michaelianblack Actually, given the corrupt election, we should have a re-vote."
Justica4all|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
morimorisdead|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
christinelu|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
christinelu|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
neilhenderson|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
neilhenderson|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
LeonidKotlyar|tass|0.5267|0.0|0.673|0.327|Legislature speaker winning presidential election in Moldovas https://t.co/US5cUbY3Uk
lawyerashley|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
PBG2017|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
sun3334|CyberkovCEO|0.0|0.0|1.0|0.0|RT @CyberkovCEO:                  !https
chulesee|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
chulesee||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
ebonieyes4u|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
dragonsandy1|realDonaldTrump|-0.8374|0.318|0.682|0.0|@realDonaldTrump @NBCNightlyNews @CNN FAKE NEWS AND PUTIN CORRUPTED OUR ELECTION! TELL THE ELECTORAL COLLEGE AND CONGRESS NO TRUMP EVER!!!!
insightspedia|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
folsomdweller2|andrewshamlet|-0.25|0.111|0.889|0.0|"RT @andrewshamlet: So while it is unclear in which direction the election will result, #socialmedia #politics #electionNight"
biggunz1965|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
biggunz1965|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
Sgym11111Greene|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
RobertDaPatriot|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
Juliacsk|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
SheriHerman10|jruha|0.0129|0.072|0.854|0.074|RT @jruha: Consider the source. CIA is master of disinformation. True that election was hacked but false that it was Russia? Cover for dome
harlan_county|ElectreIsMore|0.5542|0.0|0.796|0.204|@ElectreIsMore Still remember we had so much fun on election night here in the US.
bradisterrific|teeg_dougland|0.7237|0.0|0.748|0.252|This is a great thread by Kate and @teeg_dougland to show that it wasn't Russia that lost HRC the election https://t.co/mWE6AN3cr6
bradisterrific|twitter|0.7237|0.0|0.748|0.252|This is a great thread by Kate and @teeg_dougland to show that it wasn't Russia that lost HRC the election https://t.co/mWE6AN3cr6
LorenzoQ|randyprine|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
LorenzoQ|cnbc|-0.7905|0.333|0.558|0.11|RT @randyprine: Comey opposed outing Russians close to the election but destroying Hillary was fair game. SMH  https://t.co/qMuLvK4WEm
YellaDogTexan|aliasvaughn|-0.3597|0.102|0.898|0.0|"RT @aliasvaughn: 9. So stop trying with ""oh they just ""tried to influence"" the election"" and start realizing that what we're dealing with i"
dcapodice|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
peterjwu|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
peterjwu||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
kzootribune|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
ColiseumSewage|BenMank77|0.25|0.0|0.895|0.105|@BenMank77 @dcexaminer game-out that premise. It makes 0 sense. It would presume a predetermined election outcome counter to Dem. interests.
DianaGrannis|davebernstein|-0.4019|0.114|0.886|0.0|RT @davebernstein: Former CIA agent Robert Baer said any other country would hold a new election they found out they were hacked. (6/10)htt
TorySC|FoxNews|0.2732|0.122|0.704|0.174|"RT @FoxNews: BREAKING: Republican John Kennedy wins Louisiana runoff election for Senate seat, defeating Democrat Foster Campbell"
bchek833|summerbrennan|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
bchek833|t|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
amandar98716291|PrisonPlanet|-0.5106|0.191|0.809|0.0|"RT @PrisonPlanet: Post election riots: FAILED.Jill Stein recount: FAILED.Intimidation of EC members: FAILED.""Fake news"": FAILED.""Russia"
bryanbehar|twitter|-0.4767|0.209|0.696|0.095|We are talking about the theft of an American election by a foreign enemy. And no branch of govt willing to ensure https://t.co/vSTbm508SX
VikramSKumar|Independent|0.4404|0.0|0.828|0.172|RT @Independent: Donald Trump has thanked African Americans for not voting in the election https://t.co/uclbJZfb9r
VikramSKumar|independent|0.4404|0.0|0.828|0.172|RT @Independent: Donald Trump has thanked African Americans for not voting in the election https://t.co/uclbJZfb9r
jamesmurphypdx|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
jamesmurphypdx||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
ragwed12|Based_Gibson|-0.2732|0.179|0.722|0.099|RT @Based_Gibson: Give Obama some credit. He is reluctant to go along with the CIA/Clinton narrative that Russia hacked the election. Obama
TonyMcElhatton1|ericbolling|0.4728|0.0|0.872|0.128|RT @ericbolling: 20 business days since the Trump election. 12 new record highs in the Dow. Plus more economic opportunity here's a quick v
WalkerKaykay|ManMet80|-0.4404|0.139|0.861|0.0|RT @ManMet80: #CountryOverParty Im so old I remember when conspiring with Russia to influence election would be disqualifying and treason
FeltyKali|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
FeltyKali|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
jude_scout|austinfounde|0.0|0.0|1.0|0.0|RT @austinfounde: @SenSanders do you have nothing to say about the Russian interference in the election?
Tis4Ta|twitter|-0.4215|0.174|0.826|0.0|"Demand a new election? Why give Hillary who lost the election, she is trying anything to get a new election with https://t.co/yRjvoQhRXu"
MedievalRobots|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
MedievalRobots||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
martinitime1975|CounterMoonbat|-0.7184|0.231|0.769|0.0|RT @CounterMoonbat: If Russia hacked our election then lax cyber-security is yet another failure to add to Obama's legacy. It's a long list.
vickysue45|WeNeedTrump|-0.4522|0.129|0.871|0.0|"RT @WeNeedTrump: So the left cries about Russia allegedly interfering with our election. Yet, millions were donated to the Clinton Foundati"
igorb4662|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
politicsinred|EcuadorDeb|0.0|0.0|1.0|0.0|RT @EcuadorDeb: @Irwin_Elaine @_0HOUR1 Shows that if Putin really wanted to influence the election all he had to do was donate to the Clint
soundbites258|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
SHOPWHATUWANT2|ChristiChat|0.6249|0.0|0.796|0.204|RT @ChristiChat: During the electionit was great to see @SheriffClarke back up @realDonaldTrumpvia TV-rallies-bus tours &amp; RNCConvention#
liberalforeverX|SenSanders|0.0|0.0|1.0|0.0|@SenSanders @Missjayette Bernie Are you calling for a new election?
Ish|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Ish|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Rob_Melrose|Khanoisseur|-0.2263|0.087|0.913|0.0|RT @Khanoisseur: More new evidence that Comey tipped undecided voters toward Trump in last 2 weeks of the electionBiggest tamperer was th
rigsby_michelle|hectormorenco|0.0|0.0|1.0|0.0|RT @hectormorenco: REAL NEWS: CIA &amp; MSM Make Up False Allegations of Russian Election Tampering Without Evidencehttps://t.co/jEyE0fR09S -
SandyTomich|SenatorTomUdall|0.5267|0.067|0.714|0.219|RT @SenatorTomUdall: I will join lawmakers in both parties &amp; demand investigation of Russia's effort to influence presidential election. ht
WendySzy|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
Zhian2160|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Zhian2160||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
GarthDerby|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
GarthDerby||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
JoshuaRyanHub|YouTube|-0.5423|0.289|0.597|0.114|The Truth About Fake News | Russia Hacked U.S. Election For Donald Trump? https://t.co/jLJU6DluWP via @YouTube
JoshuaRyanHub|youtube|-0.5423|0.289|0.597|0.114|The Truth About Fake News | Russia Hacked U.S. Election For Donald Trump? https://t.co/jLJU6DluWP via @YouTube
pink_sprnva|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
salted3|_Makada_|-0.296|0.115|0.826|0.06|"RT @_Makada_: President-Elect Trump: It's ridiculous to say Russia intervened in the election, I think it's just another excuse. We had a m"
BTroyDMiller|PrisonPlanet|-0.3453|0.139|0.861|0.0|RT @PrisonPlanet: Russia interfered in the election! (no evidence).LEFT FREAKS OUT.Saudi Arabia provably bankrolled Clinton's campaign.
brenz1|CBNNews|0.0|0.0|1.0|0.0|RT @CBNNews: .@JoelCRosenberg says the mood in #Israel is upbeat after #DonaldTrump's victory in the #US presidential election. https://t.c
brenz1||0.0|0.0|1.0|0.0|RT @CBNNews: .@JoelCRosenberg says the mood in #Israel is upbeat after #DonaldTrump's victory in the #US presidential election. https://t.c
3J1963|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
xseane|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
rimaanabtawi|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
CathyLocke911|BreitbartNews|-0.1531|0.074|0.926|0.0|"RT @BreitbartNews: CORRECTION: After feedback from several Twitter folks, we now know there are NOT frequent food shortages in Ghana. https"
ElfGrove|DanielleMuscato|0.7184|0.0|0.778|0.222|"RT @DanielleMuscato: ""If Hillary Clinton won the election &amp; CIA report came out of foreign tampering, I'm sure @GOP'd be having exact same"
girls_smarter|rmasher2|-0.6486|0.227|0.773|0.0|"RT @rmasher2: If there's no constitutional mechanism to redo an election compromised by foreign interference, something's wrong with our Co"
Patta47cake|leahmcelrath|-0.3412|0.112|0.888|0.0|RT @leahmcelrath: NYTimes Editorial Board takes a stand &amp; even calls Trump out for not supporting an investigation into Russia hackinghttp
JChrisPires|brianbeutler|0.34|0.0|0.888|0.112|"RT @brianbeutler: ""Goldman Sachs has accounted for nearly a third of the Dow Jones industrial average's gains since the election. https://"
JChrisPires||0.34|0.0|0.888|0.112|"RT @brianbeutler: ""Goldman Sachs has accounted for nearly a third of the Dow Jones industrial average's gains since the election. https://"
satish_jha|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
satish_jha|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
GloriaMiele|rwindrem|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
GloriaMiele|nbcnews|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
briansonfire|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
briansonfire|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
Goodnightma|America_1st_|0.0|0.0|1.0|0.0|RT @America_1st_: BREAKING#RussianHacker was caught on camera at voting booth trying to influence election by voting for Donald J. Trum
pl8ofshrimp|MrDane1982|0.0|0.0|1.0|0.0|@MrDane1982 https://t.co/AtlfkHh7r1
pl8ofshrimp|petitions|0.0|0.0|1.0|0.0|@MrDane1982 https://t.co/AtlfkHh7r1
DeburghValerie|SarahPalinUSA|0.3254|0.131|0.657|0.211|"@SarahPalinUSA LOL   I guess you missed them messing with the election,  you r such a tool."
NijimaSan|leahmcelrath|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
NijimaSan|t|0.0|0.0|1.0|0.0|"RT @leahmcelrath: Alexandr Dugin has a Facebook page.Days after the U.S. election, he posted ""So. Washington is ours."" https://t.co/Brf1c"
LFScott57|activist360|-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
LFScott57||-0.5719|0.199|0.732|0.07|RT @activist360: Trump trashes CIA: Tries to convince his dirt dumb bigot base that Russia did not hack election to get him elected https:/
brenrey85|HuffPostPol|0.0|0.0|1.0|0.0|"Donald Trump says it is ""ridiculous"" to say Russia intervened in the election on his behalf. https://t.co/4fjQBm9JzY # via @HuffPostPol"
brenrey85|huffingtonpost|0.0|0.0|1.0|0.0|"Donald Trump says it is ""ridiculous"" to say Russia intervened in the election on his behalf. https://t.co/4fjQBm9JzY # via @HuffPostPol"
yanachoen|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
yanachoen|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
jodi_yoho|JudgeJeanine|0.0|0.0|1.0|0.0|"RT @JudgeJeanine: ""The election is over - you're either with us or against us. That is...with the U.S. or against the U.S.""-@JudgeJeanine #"
RESTORD|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
allyauriemma|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
allyauriemma|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
TxsleuthUSA|DavidAFrench|-0.3612|0.122|0.878|0.0|RT @DavidAFrench: What's the argument against a bipartisan investigation of Russian efforts to disrupt and/or influence the election? Is th
lycoris_aurea|JasonKander|-0.6597|0.213|0.787|0.0|"RT @JasonKander: If we ignore Russian espionage in our election, we embolden other foreign powers to launch similar attacks on every aspect"
Zhian2160|LindseyGrahamSC|-0.0572|0.06|0.94|0.0|"RT @LindseyGrahamSC: I'm not challenging the outcome of the election, but very concerned about Russian interference/actions at home &amp; throu"
BarryHingley|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
TroyBlayne|_HankRearden|-0.5809|0.152|0.848|0.0|"@_HankRearden @Evan_McMullin Is the CIA working with Obama to influence the election? This is the question, if so it's a high crime #MAGA"
hotmerthanyou|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
yh_boii|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Eonkidz|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
Eonkidz|t|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
ramseyellismd|VABVOX|-0.296|0.091|0.909|0.0|RT @VABVOX: 6) Trump's ties to Putin have always been suspect. Now his election's been revealed to have likely been orchestrated by a forei
LaLaLeans|intlspectator|0.3182|0.0|0.874|0.126|RT @intlspectator: Statement from prominent Republican and Democratic Senators on allegations of Russian involvement in election. https://t
LaLaLeans||0.3182|0.0|0.874|0.126|RT @intlspectator: Statement from prominent Republican and Democratic Senators on allegations of Russian involvement in election. https://t
danilo_gesmundo|danilogesmundo|0.0|0.0|1.0|0.0|Donald Trump says CIA charge Russia influenced election is 'ridiculous' - https://t.co/8XWN4z8n80 https://t.co/mhq7gfC0gx
FatAcrobat|iamaroadtrip|-0.3089|0.111|0.889|0.0|"@iamaroadtrip this account hasn't been active since 2011. It started tweeting about trump on December 3rd 2016, wel https://t.co/8E412WJOAA"
FatAcrobat|twitter|-0.3089|0.111|0.889|0.0|"@iamaroadtrip this account hasn't been active since 2011. It started tweeting about trump on December 3rd 2016, wel https://t.co/8E412WJOAA"
RevRigatone|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
GARYHARTMAN|armed-services|0.0|0.0|1.0|0.0|"McCain, Graham, Schumer, Reed Joint Statement on Reports That Russia Interfered with the 2016 Election:  https://t.co/X8iQnDWN1L"
chibi_missy|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
chibi_missy|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
christina_hikes|NewYorker|0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
christina_hikes||0.5122|0.0|0.858|0.142|"RT @NewYorker: The election of Donald Trump to the Presidency is nothing less than a tragedy for America, David Remnick writes. https://t.c"
klarson980|DavidYankovich|-0.296|0.109|0.891|0.0|RT @DavidYankovich: There is no Democrat/Republican side to the Russian influence in this election.You are either a patriot or a traitor.
therealbiostate|An0nKn0wledge|-0.6908|0.289|0.619|0.093|RT @An0nKn0wledge: Crazy Thought What If The CIA Yelled #RussiaHacking To Distract From REAL Election Fraud In Favor Hillary &amp; DHS Attempte
RobietheCat42|michaelianblack|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
RobietheCat42|twitter|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
PaulBauer21|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
tarttwit|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
steve_boyar|pgrandee10|0.0|0.0|1.0|0.0|RT @pgrandee10: @KyleNeven1 @funder Foreign involvement. The election should be invalidated. GOP corruption helped to get him elected...cou
going2left|DavidYankovich|-0.296|0.109|0.891|0.0|RT @DavidYankovich: There is no Democrat/Republican side to the Russian influence in this election.You are either a patriot or a traitor.
tekstar77|andieiamwhoiam|0.5267|0.065|0.75|0.185|"RT @andieiamwhoiam: Sorry Lefties, Russians, recounts, aliens (the extraterrestrial kind)...you will never get a new election.  Trump won."
kcimary|BreitbartNews|-0.822|0.434|0.495|0.071|RT @BreitbartNews: Why do Democrats want a war with Russia so badly? https://t.co/KfMP9vzZsu
kcimary|breitbart|-0.822|0.434|0.495|0.071|RT @BreitbartNews: Why do Democrats want a war with Russia so badly? https://t.co/KfMP9vzZsu
e_revolutionist|ImEmmaE|0.2023|0.0|0.904|0.096|RT @ImEmmaE: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/wrXVYR
e_revolutionist|t|0.2023|0.0|0.904|0.096|RT @ImEmmaE: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/wrXVYR
frankin46|frankin46|0.0|0.0|1.0|0.0|RT @frankin46: @NancyPelosi how come you guys didn't do anything before the election? Closing the barn door after the horse has gotten away
sheenA_8886|aliasvaughn|-0.2732|0.126|0.795|0.079|RT @aliasvaughn: 10. #AuditTheVote people told you straight the day after election that Russian hackers were attacking US on election night.
CarolLpr|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
CarolLpr|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
BAJVisser|nytimes|0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
BAJVisser||0.6124|0.106|0.63|0.264|RT @nytimes: A remarkable breach has emerged between Trump and intelligence agencies over claims that Russia hacked the election https://t.
crose84|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
newacademic|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
newacademic|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
folsomdweller2|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
YvonneSheffield|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
YvonneSheffield||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
hsummer|ChrisJZullo|-0.5532|0.258|0.597|0.145|RT @ChrisJZullo: Just had a dream. Republicans didn't steal the election from Al Gore. No IRAQ war or 1% tax cut. New bank regulations and
RPolsenberg|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
DebDake|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
nak006|BarkerTV|0.3182|0.0|0.916|0.084|"RT @BarkerTV: HRC: ""if we were going to push an election [in Palestine], we should have made sure that we did something to determine who wa"
postofficetruth|CNNPolitics|0.0|0.0|1.0|0.0|"RT @CNNPolitics: BREAKING: President Obama has ordered a full review into 2016 election hacking by the Russians, Lisa Monaco says https://t"
postofficetruth||0.0|0.0|1.0|0.0|"RT @CNNPolitics: BREAKING: President Obama has ordered a full review into 2016 election hacking by the Russians, Lisa Monaco says https://t"
nittmoe|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
ac_de_|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
lindadoherty4|Khanoisseur|-0.2263|0.087|0.913|0.0|RT @Khanoisseur: More new evidence that Comey tipped undecided voters toward Trump in last 2 weeks of the electionBiggest tamperer was th
dexter_zee|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
cussetabraswell|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
mattiOgreen|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
marcylauren|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
bridgeth_bro|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
bridgeth_bro|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
JustMeinMI|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
brenz1|_Makada_|-0.9081|0.383|0.617|0.0|RT @_Makada_: The same fake news media who said Iraq had weapons of mass destruction now claims Russia hacked our election. MSM are known l
CharaCarbone|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
CharaCarbone|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
AmericanSoWoke|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
rk55mk|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
FunnygirlLee|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
JosephMGindi|dailycaller|-0.3182|0.15|0.85|0.0|FBI Disagrees With CIA On Russian Influence In The Presidential Election https://t.co/FU6031FxRX via @dailycaller
JosephMGindi|dailycaller|-0.3182|0.15|0.85|0.0|FBI Disagrees With CIA On Russian Influence In The Presidential Election https://t.co/FU6031FxRX via @dailycaller
Aszneth|Bipartisan|0.0|0.0|1.0|0.0|"BREAKING: Mitch McConnell Implicated In Russia/Trump Election Meddling, FBI Inquiry https://t.co/wngmlUwSMQ via @Bipartisan Report"
Aszneth|bipartisanreport|0.0|0.0|1.0|0.0|"BREAKING: Mitch McConnell Implicated In Russia/Trump Election Meddling, FBI Inquiry https://t.co/wngmlUwSMQ via @Bipartisan Report"
SheWho__|petitions|0.0|0.0|1.0|0.0|SCOTUS: Invalidate Election Results Of 2016 - Order A New Election https://t.co/tW44ExOUxi
AlshehmaniA|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
AlshehmaniA|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
MarieMurcelle1|AnthonyTauro1|0.2003|0.167|0.625|0.208|"RT @AnthonyTauro1: @Greg_Palast Greg Palast ,crosscheck purged7.2 mil votes4 DJT, HRC won , election stolen!"
Ikipr|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Ikipr|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Granby01|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ProfChrisMJones|NickKristof|0.0|0.0|1.0|0.0|"As an academic, Trump's election was a wake-up call to me, but not for the reasons that @NickKristof seems to think. https://t.co/TYIl5P3wsZ"
ProfChrisMJones|nytimes|0.0|0.0|1.0|0.0|"As an academic, Trump's election was a wake-up call to me, but not for the reasons that @NickKristof seems to think. https://t.co/TYIl5P3wsZ"
pdcIV|BruceBartlett|0.0|0.0|1.0|0.0|"RT @BruceBartlett: The question isn't why Russia interfered in our election, the question is why did in interfere on behalf of Trump &amp; the"
Aurora_Hernandz|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
Aurora_Hernandz||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
crossfitnans|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
crossfitnans|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
randyschwart|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
ScottCross22|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
oklahomadude|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
_BuddhistPunk_|KungFunny|-0.8074|0.249|0.751|0.0|"RT @KungFunny: if russia interferred in our election, we should be investigating the hell out of it, regardess of who or what the hacked, f"
rimidott|xXSkyeCatXx|0.7184|0.0|0.684|0.316|the one good thing that came out of the election was i became friends with @xXSkyeCatXx
Connected716|summerbrennan|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
Connected716|t|0.0|0.0|1.0|0.0|"RT @summerbrennan: This is real, I checked. It's Putin's Bannon, gloating that ""Washington is ours"" after the election. https://t.co/w5w06Z"
mercedesfduran|ParkerMolloy|-0.5067|0.17|0.83|0.0|"RT @ParkerMolloy: ""patrioteagle.flag says there's a child sex pizza dungeon!""""On it!""""The CIA says Russia messed w/ the election!""Some s"
RivalThoughtsTo|DavidAFrench|0.0|0.0|1.0|0.0|@DavidAFrench You're fishing in order to overturn an election
Groovehare|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
Groovehare|washingtonpost|-0.3724|0.164|0.836|0.0|RT @washingtonpost: Trump defends his practice of not receiving a daily intelligence briefing https://t.co/w1IYcgXNPp https://t.co/49t1oYSd
crazyhorse2126|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
jjmplsmn|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
jbtcarolina|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Skrewface27|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
going2left|VABVOX|0.0|0.0|1.0|0.0|"RT @VABVOX: .@SpeakerRyan is tweeting about overturning #Obamacare, not Russian interference with our election. https://t.co/4SirvxWCKi"
going2left|twitter|0.0|0.0|1.0|0.0|"RT @VABVOX: .@SpeakerRyan is tweeting about overturning #Obamacare, not Russian interference with our election. https://t.co/4SirvxWCKi"
theSopranoist|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
theSopranoist||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
zgoelman|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
ChrisVoeller1|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
susyquu|hautedamn|-0.34|0.113|0.833|0.054|RT @hautedamn: The people who want you to believe Russia hacked the election are the same people telling you #pizzagate isn't real.
CherylDuggan1|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Mikew1767|JuddLegum|0.0|0.0|1.0|0.0|Trump adviser suggests election hacks were false flag operation by the Obama administration by @JuddLegum https://t.co/YjjsM8jTqK
Mikew1767|medium|0.0|0.0|1.0|0.0|Trump adviser suggests election hacks were false flag operation by the Obama administration by @JuddLegum https://t.co/YjjsM8jTqK
JulesMyth1970|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
juniperbreeze07|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
sgossage09|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
sgossage09||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
rwdcsw|mtracey|0.2617|0.11|0.746|0.144|"@mtracey 'We need a new election, but won't give you details, but just trust us, but don't bring up all the times we've lied &amp; manipulated.'"
MilesDon|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
MyNameIsSergius|nytopinion|0.2944|0.0|0.897|0.103|"@nytopinion So when Obama said he'd be more flexible after the election, what does that make him? https://t.co/bekdhBO7kF via @Reuters"
MyNameIsSergius|reuters|0.2944|0.0|0.897|0.103|"@nytopinion So when Obama said he'd be more flexible after the election, what does that make him? https://t.co/bekdhBO7kF via @Reuters"
IndependPress|bbc|0.0|0.0|1.0|0.0|Macedonia election: Conservatives edge ahead as votes counted - BBC News https://t.co/pdaRIFuWvj
rachie_claire|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
rachie_claire|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Txwench|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
progunz_1|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
progunz_1|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
GerardoHGarcia|JBurtonXP|-0.4019|0.124|0.876|0.0|"RT @JBurtonXP: Always remember that by ""hacked the election,"" these people mean ""released 100% authentic documents that showed real Democra"
AllDayAMazing|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
AllDayAMazing|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
SlobKebab|WalkingDead_AMC|0.4926|0.0|0.803|0.197|@WalkingDead_AMC This makes me feel better about election 2016 results ! #TheWalkingDead #reunited @AMCTalkingDead @hardwick 
billc100|kendram75|-0.4912|0.241|0.646|0.113|"RT @kendram75: Hillary Election Loss Blamed on ""Russian Hackers"" https://t.co/WylWZVbL7N obama bein the hypocrite he is!! muh russia lol"
billc100|youtube|-0.4912|0.241|0.646|0.113|"RT @kendram75: Hillary Election Loss Blamed on ""Russian Hackers"" https://t.co/WylWZVbL7N obama bein the hypocrite he is!! muh russia lol"
threespeedgirl|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
threespeedgirl|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Supertoaste|DistanceRun|0.2732|0.0|0.92|0.08|RT @DistanceRun: @politico well give him a break he's about to go down in infamy over his collusion with Putin and Comey to fix the electio
pantog|MissLizzyNJ|-0.952|0.53|0.47|0.0|"RT @MissLizzyNJ: #ImStillNotOver the fact that I lost the election because I'm a lying criminal and America hates me, so I'll blame fake ne"
daviottenheimer|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
daviottenheimer|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
ThomasBialek2|chuckwoolery|-0.4767|0.147|0.853|0.0|RT @chuckwoolery: Why are Dems crying? They handed the election to #Trump. Find out how on a new #BluntForceTruth. https://t.co/ibMBVwfms4
ThomasBialek2|bluntforcetruth|-0.4767|0.147|0.853|0.0|RT @chuckwoolery: Why are Dems crying? They handed the election to #Trump. Find out how on a new #BluntForceTruth. https://t.co/ibMBVwfms4
naveencool1998|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
Truman_Town|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
emmiehobbs0|Hispanics16|-0.5994|0.187|0.813|0.0|RT @Hispanics16: RINO War Hawks Lindsey Graham and John McCain Call for Investigation of Russia Influencing Election https://t.co/W8ZKv1uGx
emmiehobbs0|t|-0.5994|0.187|0.813|0.0|RT @Hispanics16: RINO War Hawks Lindsey Graham and John McCain Call for Investigation of Russia Influencing Election https://t.co/W8ZKv1uGx
Jimhengstenberg|RichardGrenell|0.0|0.0|1.0|0.0|"RT @RichardGrenell: Tip for @RyanLizza: If US had evidence that the Russian Government interfered with our election, we would see multiple"
mattiOgreen|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
upforhill|JoyAnnReid|0.0|0.0|1.0|0.0|"RT @JoyAnnReid: And by the way if @SenatorReid is right, and the head of the FBI stood by and let Russia meddle in our election (then did s"
sannewman|joe_smania|-0.6486|0.275|0.725|0.0|"@joe_smania I don't know. Maybe just because, post-election, anti-Trump people are ten times as paranoid and angry?"
Mother_Oya|DavidAFrench|-0.3612|0.122|0.878|0.0|RT @DavidAFrench: What's the argument against a bipartisan investigation of Russian efforts to disrupt and/or influence the election? Is th
DJT_ChosenbyGod|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
MarieMurcelle1|twitter|-0.4939|0.186|0.814|0.0|Breaking NewsPress Conference tommorow 9:30amGreg Palast-  Then meeting with DOJ about stolen electionDetails Be https://t.co/HvRZZT0wWZ
FeminismUSTD|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
FirestormOmega|KimRippere|-0.357|0.121|0.879|0.0|"RT @KimRippere: They knew abt #RussianHacking in advance, keeping it quiet=disservice. Such tainted election results not in our interest. #"
Barkforlove1|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
cheeseboot|pattonoswalt|0.4939|0.0|0.882|0.118|"RT @pattonoswalt: Seems to me, you didn't wanna talk about it before the election. Seems to me, you just turned your pretty head &amp; walked a"
MaureenCKelly|JoyAnnReid|0.0|0.0|1.0|0.0|RT @JoyAnnReid: Other than @LindseyGrahamSC is there a single principled Republican in Washigton? Russia directly intervened in our electio
Moissez1|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
llecrupnosidam|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
Chaparro916|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
vivigold197|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Tabitha__Lily|andieiamwhoiam|0.5267|0.065|0.75|0.185|"RT @andieiamwhoiam: Sorry Lefties, Russians, recounts, aliens (the extraterrestrial kind)...you will never get a new election.  Trump won."
LarryPinkerton|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
kazpaul49|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
kazpaul49||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
micahsgrrl|DailyNewsBin|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
micahsgrrl|palmerreport|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
SFinEville|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
SFinEville|esquire|-0.2057|0.131|0.869|0.0|RT @esquire: Russia's interference in this election should not be a surprise https://t.co/Ue0oToG8rh https://t.co/ysGRqJcN8s
3Panda3|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
emilyfearnow|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
mommyofboys4|MMFlint|0.8689|0.077|0.568|0.355|RT @MMFlint: The CIA has determined Russia hacked into our election to help elect Donald J. Trump. Now Trump names Putin best friend as OUR
aprov2480|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
janiceponchak|powerlineblog|-0.5319|0.462|0.538|0.0|"People, emails were HACKED  https://t.co/obGbUbU2gl"
BrendaFiles2|mtracey|-0.7003|0.315|0.58|0.105|RT @mtracey: I assumed the crackpot Russia hysteria would subside somewhat after the election. I was wrong. People have truly gone insane.
FanciFlautist|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
Cindyg1948Cindy|jasonmurphynat1|0.0|0.0|1.0|0.0|"RT @jasonmurphynat1: @JohnTDolan @jojoh888 Yet, Obama interfered in Israel's election and McCain did NOT call for an investigation."
msjbe20a|StopTheSpeaker|0.6705|0.0|0.776|0.224|"RT @StopTheSpeaker: Paul Ryan at odds with the GOP who oversee intelligence, Pentagon and Homeland Security - Russia meddled in election ht"
aliasvaughn|twitter|-0.2263|0.095|0.905|0.0|This petition demanding a new election with paper ballots needs 100k signatures before EC votes. If you can spare a https://t.co/bCxNtLzp0A
vlassover|nytimesworld|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
vlassover|nytimes|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
sheenA_8886|aliasvaughn|-0.3597|0.102|0.898|0.0|"RT @aliasvaughn: 9. So stop trying with ""oh they just ""tried to influence"" the election"" and start realizing that what we're dealing with i"
GNSNick|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
MooreFay|thehill|0.0|0.0|1.0|0.0|FBI breaks with CIA on Russia interference in U.S. election https://t.co/BbW9dMPtot
hatekillshate|leahmcelrath|0.5584|0.0|0.796|0.204|RT @leahmcelrath: Watergate seems like such an minor almost innocent bit of subterfuge compared to what's happened in this election.
BDR121068|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
BDR121068|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
mtighe15|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
mtighe15|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
bagglo|WeAreAlreadyGr1|-0.9106|0.404|0.596|0.0|"RT @WeAreAlreadyGr1: You're a stooge amongst many stooges. Not pissed about election, just LOATHE assho*les, thugs, &amp; liars. Unlike $, your"
2ALAW|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
MuathAyesh|BrookingsInst|0.0|0.0|1.0|0.0|RT @BrookingsInst: 46% of Americans think Obama should take action on Israel-Palestine before leaving office https://t.co/pr01irnpBj https:
MuathAyesh|brookings|0.0|0.0|1.0|0.0|RT @BrookingsInst: 46% of Americans think Obama should take action on Israel-Palestine before leaving office https://t.co/pr01irnpBj https:
therealbiostate|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
therealbiostate|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
drjanet|DeanJulie|-0.2247|0.19|0.645|0.164|RT @DeanJulie: You know if HRC won &amp; CIA said Russia helped you'd be losing your fucking shit right now. This is a coup = NOT okay. https:/
drjanet||-0.2247|0.19|0.645|0.164|RT @DeanJulie: You know if HRC won &amp; CIA said Russia helped you'd be losing your fucking shit right now. This is a coup = NOT okay. https:/
KirstinElaine1|DrJillStein|0.0|0.0|1.0|0.0|"RT @DrJillStein: We expect bank tellers to double-check money before handing it to us. Let's double-check election results, too. #Recount20"
_flanders|ZaibatsuNews|0.2023|0.0|0.904|0.096|RT @ZaibatsuNews: WATCH: Chuck Todd hammers Reince Priebus over refusal to admit Russians might have influenced election https://t.co/ZuFWJ
_flanders|t|0.2023|0.0|0.904|0.096|RT @ZaibatsuNews: WATCH: Chuck Todd hammers Reince Priebus over refusal to admit Russians might have influenced election https://t.co/ZuFWJ
Ksodeeya|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
Ksodeeya|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
tomatosalad64|SenatorTomUdall|0.5267|0.067|0.714|0.219|RT @SenatorTomUdall: I will join lawmakers in both parties &amp; demand investigation of Russia's effort to influence presidential election. ht
Nicole__MarieeG|cctvnews|-0.3612|0.135|0.865|0.0|RT @cctvnews: Donald Trump: CIA assessment of Russian interference in US election ridiculous. Follow us for updates.
jwdsfca13|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
jwdsfca13||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
HonorFounders|slate|-0.34|0.156|0.844|0.0|Key senators: Reports of Russian election meddling should alarm every American. https://t.co/pD3lSgXg9e via @slate
HonorFounders|slate|-0.34|0.156|0.844|0.0|Key senators: Reports of Russian election meddling should alarm every American. https://t.co/pD3lSgXg9e via @slate
ggrushko|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
tahino1|PuestoLoco|0.0|0.0|1.0|0.0|RT @PuestoLoco: .@BillClinton spits it out: Putins boy - @FBIs James Comey is a traitor.https://t.co/DjRK7rYsoJ https://t.co/hJ5KOXMLGM
tahino1|twitter|0.0|0.0|1.0|0.0|RT @PuestoLoco: .@BillClinton spits it out: Putins boy - @FBIs James Comey is a traitor.https://t.co/DjRK7rYsoJ https://t.co/hJ5KOXMLGM
ItsMeCathi|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
Juliacsk|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
hollowman777|_HankRearden|-0.8176|0.309|0.691|0.0|@_HankRearden @TroyBlayne His candidate of choice lost (even with his fake Presidency bid) and now his butt hurts and wants a 2nd election.
HeidiJaster|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
MoChroi1965|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
MoChroi1965|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
malakim2099|ashleylynch|-0.4404|0.127|0.873|0.0|@ashleylynch I've been linking the end of that movie too much as a reaction to events after the US Election Day. :(
Anyshka|HRCNJVolunteers|-0.4215|0.135|0.865|0.0|RT @HRCNJVolunteers: @GoddessKerriLyn @srauer20 Trump disqualified self. Election had 2 candidates. 1's out. By default it's HRC in now. #S
bigfortiesfan|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
Pennie_Bennie|girlsreallyrule|0.4215|0.056|0.821|0.123|"RT @girlsreallyrule: Trump colluded with #RussianHackers to rig a free election all under the watch of Comey, the HEAD OF THE FBI and HE DI"
throbbin_willy|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Perezdog968Mike|ejenk|0.7906|0.0|0.696|0.304|RT @ejenk: I saw a video of Russians cheering on the rooftops in New Jersey when Trump won the election.
leftoftheright|BryanDawsonUSA|-0.3612|0.135|0.865|0.0|RT @BryanDawsonUSA: GOP Congress:Hearings on #Benghazi witch hunt: 33Hearings on real Russian interference in US election: 0#russianha
Th2shay|SheriHerman10|-0.4939|0.198|0.802|0.0|@SheriHerman10 The CIA are mad at Comey's FBI letters. CIA on Clinton's team.Comey https://t.co/59U0c8WK5l
Th2shay|independent|-0.4939|0.198|0.802|0.0|@SheriHerman10 The CIA are mad at Comey's FBI letters. CIA on Clinton's team.Comey https://t.co/59U0c8WK5l
MarcIntheOC|trex9123|-0.5423|0.191|0.809|0.0|RT @trex9123: @NPR @jasunmark There need to be mass resignations by editors/producers at all major media outlets who mostly ignored story d
7bugglettes|emigre80|-0.3802|0.217|0.662|0.121|"RT @emigre80: Both Trump and Sanders were delighted to cry ""rigged election!"" when they ran against Clinton.Now that there's evidence? *C"
theirishdiet|Shakestweetz|0.7165|0.105|0.64|0.255|RT @Shakestweetz: It's quite an amazing sight watching the party who sainted Ronald Reagan show an aggressive indifference to Russian inter
PoliticsUSTD|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Juliette_Rulz|KanamynLogic|0.4703|0.0|0.765|0.235|"RT @KanamynLogic: @RT_com @SputnikInt campaigning is not quite election tampering, lol"
CindyRae1960|AlexMohajer|0.5511|0.0|0.754|0.246|"RT @AlexMohajer: ""The truth? @HillaryClinton did not lose the 2016 presidential election. We did."" @HuffingtonPost https://t.co/uGErzEPz9T"
CindyRae1960|huffingtonpost|0.5511|0.0|0.754|0.246|"RT @AlexMohajer: ""The truth? @HillaryClinton did not lose the 2016 presidential election. We did."" @HuffingtonPost https://t.co/uGErzEPz9T"
SrayOrman|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
SrayOrman|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
crossfitnans|politico|0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
crossfitnans||0.4588|0.195|0.496|0.309|RT @politico: Trump calls intelligence reports of election meddling ridiculous. But prominent senators from both parties disagree https://t
vesperview|HillaryClinton|-0.7717|0.339|0.661|0.0|"First @HillaryClinton lost because of Russia, then she lost because of ""fake news"", now it's the FBI. https://t.co/JGouTAx5UF"
vesperview|thehill|-0.7717|0.339|0.661|0.0|"First @HillaryClinton lost because of Russia, then she lost because of ""fake news"", now it's the FBI. https://t.co/JGouTAx5UF"
TheHardMan21|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
heather2kin|PrisonPlanet|-0.2003|0.116|0.797|0.087|"@PrisonPlanet HR Clinton! 1: payback for her interference in their election 2. She's weak &amp; can be bought, Putin could easily count on doing"
JoferJoseph|Khanoisseur|-0.2263|0.087|0.913|0.0|RT @Khanoisseur: More new evidence that Comey tipped undecided voters toward Trump in last 2 weeks of the electionBiggest tamperer was th
_RaulRevere|mitchellvii|-0.7351|0.22|0.78|0.0|RT @mitchellvii: I don't get it.  The Media is using the same attacks against Trump that failed during the election.  They need to hire bet
Chrismf6|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
Chrismf6|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
MeredithMarsha1|TexIrvin|0.4624|0.122|0.636|0.242|@TexIrvin I hope the DNC elects him--the gift that keeps on giving-to Conservatives--they'll never win another National election or States!
tlduke_rph|NotJoshEarnest|0.471|0.0|0.861|0.139|"RT @NotJoshEarnest: Listen up folks! Just because we lie about everything, doesn't mean we're lying about Russia hacking the election."
merikab|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
lasershow109|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
lasershow109|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
maxasteele|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
DavidAWeinberg|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
DavidAWeinberg||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
airforce2100|realDonaldTrump|0.6249|0.0|0.83|0.17|"RT @realDonaldTrump: I spent Friday campaigning with John Kennedy, of the Great State of Louisiana, for the U.S.Senate. The election is ove"
PSBbazmalea|YouTube|0.0|0.0|1.0|0.0|HAITI NEWS ELECTION 2016 GADE KI SA KI RIVE Arisitid: https://t.co/a6I4lHdJCk via @YouTube
PSBbazmalea|youtube|0.0|0.0|1.0|0.0|HAITI NEWS ELECTION 2016 GADE KI SA KI RIVE Arisitid: https://t.co/a6I4lHdJCk via @YouTube
BrianCarroll89|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
BrianCarroll89|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
UWantMyVote_Why|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
UWantMyVote_Why|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
jumpouttheboat|occupydemocrats|0.0|0.0|1.0|0.0|Of course. https://t.co/3i1N3bunus
politicsinred|Irwin_Elaine|0.0|0.0|1.0|0.0|RT @Irwin_Elaine: @_0HOUR1 Here's a list of all the Foreign Governments who interfered in the last Pres election. I mean... donated to the
lindadoherty4|Khanoisseur|0.0|0.0|1.0|0.0|"RT @Khanoisseur: Not only did Trump ask Russia to hack a political rival, he took millions from them before the election @1liners https://t"
lindadoherty4||0.0|0.0|1.0|0.0|"RT @Khanoisseur: Not only did Trump ask Russia to hack a political rival, he took millions from them before the election @1liners https://t"
Teamnguns|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
OWSTimes|google|0.0|0.0|1.0|0.0|Hillary Was More Abigail Adams than Eleanor Roosevelt. That May Have Cost Her the Election. https://t.co/sAffiiSiKv  - #ows
LindaMarkss|DavidYankovich|-0.296|0.109|0.891|0.0|RT @DavidYankovich: There is no Democrat/Republican side to the Russian influence in this election.You are either a patriot or a traitor.
smell3roses|ZaibatsuNews|0.2023|0.0|0.904|0.096|RT @ZaibatsuNews: WATCH: Chuck Todd hammers Reince Priebus over refusal to admit Russians might have influenced election https://t.co/ZuFWJ
smell3roses|t|0.2023|0.0|0.904|0.096|RT @ZaibatsuNews: WATCH: Chuck Todd hammers Reince Priebus over refusal to admit Russians might have influenced election https://t.co/ZuFWJ
WillPinkston|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
cacisa2j|michaelianblack|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
cacisa2j|twitter|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
JillStorey2020|GlenFrost|0.8225|0.0|0.714|0.286|RT @GlenFrost: Why did Trump win? Richard Wolff explains before the US election why Trump was going to win https://t.co/qUasgLCzon (note; 1
JillStorey2020|youtube|0.8225|0.0|0.714|0.286|RT @GlenFrost: Why did Trump win? Richard Wolff explains before the US election why Trump was going to win https://t.co/qUasgLCzon (note; 1
BITW140|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
BITW140|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Douga536|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
ScotClimate|medium|0.0|0.0|1.0|0.0|ClimateProgress:Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/apAc3sr95v
matthew1nelson1|JIanoale|0.3182|0.0|0.901|0.099|@JIanoale the election is over and he's not president yet so he doesn't need my votes and obama can still pardon Hillary
preachingterp|CNN|-0.5106|0.292|0.708|0.0|Where's the outrage over the Russia hack? @CNN https://t.co/uqyGzy3qO1
preachingterp|cnn|-0.5106|0.292|0.708|0.0|Where's the outrage over the Russia hack? @CNN https://t.co/uqyGzy3qO1
vancitydan|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
vancitydan|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
PlantsLoveCO2|medium|0.0|0.0|1.0|0.0|ClimateProgress:Trump adviser suggests election hacks were false flag operation by the Obama administration https://t.co/7oQlLfXvDJ
mercedesfduran|mizmaxgordon|0.0|0.0|1.0|0.0|RT @mizmaxgordon: Still think Russia had nothing to do with rigging the election? Read this entire thread. #WeveBeenPwned #IllegitimateElec
allisonpowers13|AliciaDede|0.0|0.0|1.0|0.0|RT @AliciaDede: Foreign Governments who donated for Hillary's Foundation did not interfere with the election? https://t.co/JjR9yNaVNQ
allisonpowers13|twitter|0.0|0.0|1.0|0.0|RT @AliciaDede: Foreign Governments who donated for Hillary's Foundation did not interfere with the election? https://t.co/JjR9yNaVNQ
575haiku|GaryStLawrence|-0.6249|0.221|0.779|0.0|RT @GaryStLawrence: Literally EVERYONE who knew about or participated in #Russia's manipulation of our #election must be tried for treason.
CllrBSilvester|ericbolling|0.4728|0.0|0.872|0.128|RT @ericbolling: 20 business days since the Trump election. 12 new record highs in the Dow. Plus more economic opportunity here's a quick v
TroyalBrown|twitter|0.7269|0.0|0.736|0.264|"I predicted 6 months ago that Trump would win.  Not sure how I knew, I just did. I also predicted on election night https://t.co/sHERekALum"
vquagliana|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
vquagliana|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
msjbe20a|DailyNewsBin|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
msjbe20a|palmerreport|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
gruesomegull|twitter|0.4238|0.122|0.653|0.224|"Never have so many friends, allies &amp; American citizens felt so uneasy by a #election With the popular vote at 2 1/2 https://t.co/KhisrhvG50"
OWNYOMAMA|Evasabe|-0.4717|0.339|0.661|0.0|@Evasabe But she didn't win the election
shortyd1717|blaubok|0.47|0.096|0.652|0.252|RT @blaubok: When her election was 98% certain - Hillary assured Trump - the election isn't riggedWhen she lost - the election was rigged
Marie____Taylor|ndtv|0.0|0.0|1.0|0.0|Donald Trump On Russia Meddling In US Election: 'I Don't Believe It' https://t.co/ndlNMooQyz
lowki|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
lowki|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
HougenJ|sjredmond|-0.7003|0.453|0.547|0.0|"@sjredmond @Amaliada Shit, was the election about TV critics?"
celticroot|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Sailfish157|mhmck|0.0|0.0|1.0|0.0|"RT @mhmck: Rerun the election. Paper ballots. Two names: Clinton, Trump. International observers by the tens of thousands. Ukraine did it."
Vote_American|thehill|0.0|0.0|1.0|0.0|"@thehill Comey's letter didn't cost Hillary the Election, Hillary cost Hillary the Election."
Tull007|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
hatrok81|fxnopinion|0.1027|0.082|0.821|0.097|"RT @fxnopinion: Last night on ""Justice,"" Judge Jeanine Pirro had stark words for those who refuse to accept the results of the 2016 preside"
flulrich|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
flulrich|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Marie____Taylor|SuryaRay|0.0|0.0|1.0|0.0|#Indian #SuryaRay Donald Trump On Russia Meddling In US Election: 'I Don't Believe It': https://t.co/lf2qB1gaNn #Indian @SuryaRay
Marie____Taylor|ndtv|0.0|0.0|1.0|0.0|#Indian #SuryaRay Donald Trump On Russia Meddling In US Election: 'I Don't Believe It': https://t.co/lf2qB1gaNn #Indian @SuryaRay
PrettyBeaches|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
PrettyBeaches||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
RobertH01920864|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
RobertH01920864|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
Newyorker2212|twitter|0.3612|0.0|0.889|0.111|Feds found the evidence of hacking.  RNC kept it hidden just like the Keir the Russian influence in election hidden https://t.co/W1rshdaJT0
JunaidNoorCPA|sarahkendzior|0.2023|0.0|0.893|0.107|"RT @sarahkendzior: Important post on Trump, Jared Kushner, data collection, and the election #Resist https://t.co/UJkJlhEtJW https://t.co/Q"
JunaidNoorCPA|m|0.2023|0.0|0.893|0.107|"RT @sarahkendzior: Important post on Trump, Jared Kushner, data collection, and the election #Resist https://t.co/UJkJlhEtJW https://t.co/Q"
beckypsowers|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
Olegnad_Nosaj|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Olegnad_Nosaj||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
scutify|scutify|0.0|0.0|1.0|0.0|3 China Stocks to Buy Before They Make a BIG Comeback https://t.co/S8TRyb25Kw $BIDU $BABA $MPEL $AMZN $TSLA $GOOG https://t.co/pKAwIgkj2h
VincentTaddei|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
maureenking79|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
maureenking79|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
dorbar|theguardian|0.0|0.0|1.0|0.0|The only transparent thing about Obama's admin is their endless efforts to over-turn democratic elections results!https://t.co/gR2p6TRFew
kppwrites|BruceBartlett|0.0|0.0|1.0|0.0|"RT @BruceBartlett: The question isn't why Russia interfered in our election, the question is why did in interfere on behalf of Trump &amp; the"
peterb442|peddoc63|0.0|0.0|1.0|0.0|RT @peddoc63: Here's a list of foreign governments that interfered with presidential election....oops I meant donated to Clinton Foundation
Kam_Holt|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Kam_Holt||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
j_danielo|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
KatrinaGrau|NCCollegians|-0.7531|0.33|0.548|0.122|RT @NCCollegians: Liberals before the election: Wow Trump is a moron. Voter fraud is just a myth. Liberals after the election: RIGGED ELE
makledes|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
makledes|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
NoGunsNoGulag|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
NoGunsNoGulag|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
ItsSeanRoach|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
raghask|girishalva|-0.1351|0.102|0.816|0.082|"RT @girishalva: In 1996,Rajinikanth said ""If Jaya is voted back 2 power, even God can't save TN"". Was it the reason for her defeat?https:/"
raghask||-0.1351|0.102|0.816|0.082|"RT @girishalva: In 1996,Rajinikanth said ""If Jaya is voted back 2 power, even God can't save TN"". Was it the reason for her defeat?https:/"
anthonytshering|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
anthonytshering||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
paul_carilli|Politikath|0.0|0.0|1.0|0.0|RT @Politikath: Ex-CIA operative: We may need a new vote @CNNPolitics https://t.co/bPZ4kcxUjn
paul_carilli|edition|0.0|0.0|1.0|0.0|RT @Politikath: Ex-CIA operative: We may need a new vote @CNNPolitics https://t.co/bPZ4kcxUjn
Devendra2555|PathiShashidhar|0.5106|0.0|0.845|0.155|RT @PathiShashidhar: @timesnow Madam #Mamata if u hv confidence y don't u dissolve ur assembly and go for election in ur State.
vquagliana|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
vquagliana|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
TeamSheaPorter|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
maganti_rk|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
DMMadora|wendyvoss|0.0|0.0|1.0|0.0|RT @wendyvoss: Immediate Attention! https://t.co/xQoUl0lu7F
DMMadora|infowars|0.0|0.0|1.0|0.0|RT @wendyvoss: Immediate Attention! https://t.co/xQoUl0lu7F
SavvDaddy|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
SavvDaddy|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
IsaacBloomberg|mat_johnson|0.4404|0.0|0.861|0.139|@mat_johnson @Bencjacobs I'll do you one better. The whole election was a false false flag operation by the Bush Administration.
The_A_Prentice|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
The_A_Prentice|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
lang3rsh|RogersParkMan|-0.3818|0.11|0.89|0.0|"RT @RogersParkMan: Hey @fakedansavage , think R's would be upset if Russians are found to have tampered with the R Primaries, not just the"
leigh_marthe|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
leigh_marthe|t|0.0|0.0|1.0|0.0|RT @wikileaks: Former UK Ambassador Craig Murray on recent anonymous CIA claims about alleged US election related sources https://t.co/LcTD
ChrisGaryL|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: CNN: Obama orders report into WikiLeaks timed for release just prior to Trump presidency https://t.co/YZNpSht3tjhttps://t.
ChrisGaryL|t|0.0|0.0|1.0|0.0|RT @wikileaks: CNN: Obama orders report into WikiLeaks timed for release just prior to Trump presidency https://t.co/YZNpSht3tjhttps://t.
zonesergio1|claudiawrites|0.2187|0.109|0.743|0.147|RT @claudiawrites: Don't betray those who gave their lives fighting for their country. Investigate Russian ties to election. #CountryOverPa
OLochlainn|RealAlexJones|-0.7865|0.348|0.652|0.0|RT @RealAlexJones: #CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia - https://t.co/eXe3mPaIEG #infowars
OLochlainn|youtube|-0.7865|0.348|0.652|0.0|RT @RealAlexJones: #CIA Election Report Is FAKE NEWS To Attack Trump &amp; Russia - https://t.co/eXe3mPaIEG #infowars
87bladesmom|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
javie26|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
cussetabraswell|Khanoisseur|0.0|0.0|1.0|0.0|"RT @Khanoisseur: Not only did Trump ask Russia to hack a political rival, he took millions from them before the election @1liners https://t"
cussetabraswell||0.0|0.0|1.0|0.0|"RT @Khanoisseur: Not only did Trump ask Russia to hack a political rival, he took millions from them before the election @1liners https://t"
EllyHuy|youtube|-0.5473|0.202|0.798|0.0|"HEATED Debate | Reince Priebus DENIES CIA Evidence of Election HACKS, ""You Can't Prove ANYTHING"" https://t.co/BfHv1gQhtH"
juannec|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
Simplysimon818|MaxSteel747|-0.6908|0.231|0.769|0.0|RT @MaxSteel747: Democrats Are Using the Same Corrupt Political System to Steal the Presidency From Trump &amp; Claim Russians Rigged Election~
marcatcar|neilpX|-0.5423|0.17|0.83|0.0|"RT @neilpX: If McCain and Graham are able to expose the treason promulgated in the election, they will deserve to be heralded as American h"
idle_prattle|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
alicia3281|robreiner|0.0|0.0|1.0|0.0|"RT @robreiner: Teapot Dome,Watergate,Iran-Contra are quaint compared to Russian gov. in league with Trump to influence US election. Crimina"
jaded_gal05|EdWorthy10|0.4265|0.0|0.898|0.102|"RT @EdWorthy10: The Electoral College Vote on Dec 19th is still the MOST important event since the election. To get to Jan 20th, we must ge"
sabrinaabv|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
PrettyBeaches|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
Amy____Jones|ndtv|0.0|0.0|1.0|0.0|Donald Trump On Russia Meddling In US Election: 'I Don't Believe It' https://t.co/U4HRMx94lz
AspiringThrawn|EscapeVelo|-0.3182|0.113|0.887|0.0|RT @EscapeVelo: The FBI leaked that #GamerGate was a Russian psyops operation designed to influence the 2016 Presidential Election. #Stop
pinklady404|kamrananwar1973|-0.6679|0.199|0.801|0.0|RT @kamrananwar1973: @Headerop1 @markoff @DailyNewsBin Then we deserve a do over!!!  Too much shit Interfered with this election and a PIG
JamesTKingP1|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
JamesTKingP1||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Cindyg1948Cindy|LibertyFolders|-0.5267|0.167|0.833|0.0|RT @LibertyFolders: Remember: Obama the hypocrite interfered in Israel's elections but he has balls 2 criticize Russia 4 supposedly interfe
EDee_1|_Makada_|0.0431|0.113|0.768|0.119|"RT @_Makada_: Obama ordered intelligence agencies to investigate Russian interference in election with NO PROOF, by doing this he is the on"
MichaelRayAdam2|NotJoshEarnest|-0.4738|0.206|0.702|0.092|"RT @NotJoshEarnest: Remember when not accepting election results was a danger to the democracy? Seems like it was last month. Oh wait, it w"
Amy____Jones|ndtv|0.0|0.0|1.0|0.0|Donald Trump On Russia Meddling In US Election: 'I Don't Believe It' https://t.co/dvC17BxJoF
justclay12|JoyAnnReid|0.4404|0.0|0.873|0.127|"RT @JoyAnnReid: Baer makes a good point: if we had been caught interfering in a foreign country's election, they would redo their election."
JaiHIndtweets|jomalhotra|0.7548|0.0|0.682|0.318|RT @jomalhotra: @manupubby_ET @manoharparrikar The Goa election campaign is more important than celebrating Navy Day by the Defence Ministe
Judigal|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
arachnea|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
arachnea||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
hello_jaime|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
RobotDeathSquad|ParkerMolloy|-0.5067|0.17|0.83|0.0|"RT @ParkerMolloy: ""patrioteagle.flag says there's a child sex pizza dungeon!""""On it!""""The CIA says Russia messed w/ the election!""Some s"
DpeltoD|ProgressiveMass|0.0|0.0|1.0|0.0|@ProgressiveMass any upcoming meetings in Boston area? Been quiet since election
blaha_b|emigre80|-0.3802|0.217|0.662|0.121|"RT @emigre80: Both Trump and Sanders were delighted to cry ""rigged election!"" when they ran against Clinton.Now that there's evidence? *C"
paul_daytripper|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Marie_Al_Marie|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
pnr9|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: Heres a list of the governments that tried to influence our election (donated to the Clinton foundation). None of thes
triplesss1001|kurteichenwald|0.0|0.0|1.0|0.0|RT @kurteichenwald: @thedailybeast Bernstein also said Comey wouldn't have announced pre-election unless something major. Woodward said ema
UNKLE_PAULEE|YouTube|-0.5859|0.213|0.787|0.0|"[40] Election Recount Shows Fraud, Veterans Stand w/ Standing Rock, &amp; De... https://t.co/J3ri7UwqH7 via @YouTube"
UNKLE_PAULEE|youtube|-0.5859|0.213|0.787|0.0|"[40] Election Recount Shows Fraud, Veterans Stand w/ Standing Rock, &amp; De... https://t.co/J3ri7UwqH7 via @YouTube"
cissy_Ike|d_fucile|-0.5449|0.133|0.867|0.0|RT @d_fucile: THERE'S NO NEW ELECTION!  THE RUSSIANS DIDN'T HACK! ONE MAN WHO WAS INVOLVED WITH ASSANGE ALREADY SAID IT WAS NOT RUSSIANS AS
mpostles|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
BigMouth1122|An0nKn0wledge|-0.6739|0.171|0.829|0.0|RT @An0nKn0wledge: THERE IS MORE EVIDENCE OF ALIENS EXISTING THEN THE RUSSIANS HACKING THE ELECTION.. BTW THE ELECTION FRAUD SO FAR ALL IN
vchartier2902|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
c_greggain|RichardGrenell|0.0|0.0|1.0|0.0|"RT @RichardGrenell: Tip for @RyanLizza: If US had evidence that the Russian Government interfered with our election, we would see multiple"
MARAUDER78|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
MARAUDER78|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
wendybyrdm|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
wendybyrdm|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
ZNittmo|MMFlint|0.8689|0.077|0.568|0.355|RT @MMFlint: The CIA has determined Russia hacked into our election to help elect Donald J. Trump. Now Trump names Putin best friend as OUR
ptrmsk|historyinflicks|-0.3612|0.106|0.894|0.0|RT @historyinflicks: Trump in Nov: the election could be rigged. i might not concede.Dems in Dec: change dot org petition asking the Deep
bannerite|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
bannerite||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
mrgasmaskman|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
mrgasmaskman|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
dah1776|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
flintr|SenatorTomUdall|0.5267|0.067|0.714|0.219|RT @SenatorTomUdall: I will join lawmakers in both parties &amp; demand investigation of Russia's effort to influence presidential election. ht
LindaMadison10|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
LindaMadison10|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
graybruce|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
graybruce||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
DMMadora|FoxNewsSunday|0.8625|0.0|0.676|0.324|RT @FoxNewsSunday: We hope you enjoyed the show today w/ President-elect Trump as he spoke in his first Sunday show interview since winning
llsmith2449|blogbooktours|-0.5904|0.193|0.807|0.0|@blogbooktours: How Russia Pulled Off the Biggest Election Hack in U.S. History https://t.co/f3oowfts9b via @Esquire FAKE NEWS
llsmith2449|esquire|-0.5904|0.193|0.807|0.0|@blogbooktours: How Russia Pulled Off the Biggest Election Hack in U.S. History https://t.co/f3oowfts9b via @Esquire FAKE NEWS
ProudDemocrat1|kurteichenwald|0.0|0.0|1.0|0.0|"RT @kurteichenwald: Also, there must be investigation of Comey @FBI. That he could know this &amp; decide to break all history to interfere w/"
srikki03|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
yunibuny1|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
morphsintowomen|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
tylr|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
tylr|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
bamilekeeavon|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
bamilekeeavon|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
wandsci|BrendanNyhan|-0.4659|0.169|0.787|0.043|"RT @BrendanNyhan: Seeing people dismiss as silly conspiracy talk, but far more serious. Potential Dep SOS suggesting Obama used IC in a dom"
Amatodeb|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
paintedparrot|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
BayouWho|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
_sean_casey|MaydnUSA|-0.4019|0.119|0.881|0.0|"RT @MaydnUSA: When Sony was hacked, the FBI immediately produced evidence. Anyone seen any actual evidence of election hack by Russia?Did"
tab24759|SonofLiberty357|-0.5267|0.152|0.848|0.0|"RT @SonofLiberty357: This is what's being called 'hacking, influencing election."" Somebody leaking emails that show the Dems to be lying, c"
DKshad0w|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
DKshad0w|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
zackmomma|ImEmmaE|0.2023|0.0|0.904|0.096|RT @ImEmmaE: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/wrXVYR
zackmomma|t|0.2023|0.0|0.904|0.096|RT @ImEmmaE: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/wrXVYR
jenfries|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
marypmadigan|foreignpolicy|0.0|0.0|1.0|0.0|It Was a Corruption Election. Its Time We Realized It. https://t.co/zQt1vpzjpi
YeeunMin1|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
WestieGal|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
RtmTweets|PolitixGal|-0.5043|0.183|0.817|0.0|RT @PolitixGal: Continued MSM claim that Russian leaks lost Clinton the election while still never acknowledging the truth the leaks reveal
TVNewsWatchDog|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
TVNewsWatchDog|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
puhi8251|phil200269|0.0|0.0|1.0|0.0|RT @phil200269: What if the election hadn't been hacked?What if Hillary hadn't stole the nomination?What if Obama hadn't given rise to
tim6731|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
tim6731||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Chris_Ledbetter|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
pwykoff|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Jojo_Lovejoy|swin24|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
Jojo_Lovejoy|thedailybeast|0.3612|0.0|0.865|0.135|"RT @swin24: like, Trump publicly did this, actually: ""Russia, if you're listening"" he said @ a rally https://t.co/u8yujY22EM https://t.co"
ge2229617|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
nancy875|eileendefreest|-0.4588|0.143|0.857|0.0|RT @eileendefreest: Mitch McConnell knew about #RussianHacking in Oct. and threatened Obama w/being partisan if data released to American v
TaKingOfAwkward|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
TaKingOfAwkward|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
duhgurlz|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
bloggoneit|WalshFreedom|0.0|0.0|1.0|0.0|RT @WalshFreedom: .@SpeakerRyan refuses to call for an investigation into Russia meddling in the election.Coward.https://t.co/hpS8ApqMfq
Konamali1|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
starknightz|twitter|-0.6486|0.29|0.71|0.0|Reince Priebus Battles NBCs Chuck Todd on Russian Election Hacking  Chuck This Is Insane https://t.co/hLEUn2G2jj
KB24xJG24|VeganLoveTeach|0.128|0.104|0.769|0.127|"RT @VeganLoveTeach: @AlexMohajer @HillaryClinton If you take CA out, she loses popular vote.  California shouldn't decide the election.  Th"
leeromney|palmerreport|-0.4215|0.128|0.872|0.0|Fifty-nine percent of the vote counting machines in Detroit -- Michigans biggest city -- all broke on Election Day. https://t.co/lJ6EQ7VndM
Minerva452010|MarkYoungTruth|-0.4976|0.295|0.58|0.125|@MarkYoungTruth @Talk2Rusty So called tolerant liberals who protest and riot after the election result.
mariespearsai|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
PollySimson|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
AppellateJunkie|lawfareblog|-0.5423|0.36|0.64|0.0|Lawfareblog's take--it's critical to respond to Russia's election aggression: https://t.co/ar7K1ecYH8
ProvaxShill|themattmcd|0.0|0.0|1.0|0.0|RT @themattmcd: Here is Mitch McConnell's office number:202-224-2541Call and ask why he kept us in the dark about foreign interference
TheborderIzsafe|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
TheborderIzsafe|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
BossClaw|JBurtonXP|-0.4019|0.124|0.876|0.0|"RT @JBurtonXP: Always remember that by ""hacked the election,"" these people mean ""released 100% authentic documents that showed real Democra"
amag88|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
D_Graettinger|PolitiFact|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
D_Graettinger|t|0.1027|0.101|0.78|0.119|RT @PolitiFact: NEW: Priebus says there's no clear report on Russia trying to shape US election. False. @MeetThePress https://t.co/YbOVAjVb
2ALAW|CarmineZozzora|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
2ALAW|t|0.2462|0.094|0.77|0.136|"RT @CarmineZozzora: Oct 31, 2016: FBI sees no clear link to Russia:https://t.co/L4av41NW2aPost Nov 8th: It was Russia! Russia did it! C"
tootropic|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
tootropic|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
rigsby_michelle|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
DKWilson56|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
janefc3|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
scrubbyscum999|JBurtonXP|0.6597|0.0|0.779|0.221|"RT @JBurtonXP: If Russia wanted to influence the election, they should've just donated millions to Hillary like all the respectable foreign"
DellaCooper3|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
DellaCooper3||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
BelisaDavis|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
r1965rainey|NotJoshEarnest|0.471|0.0|0.861|0.139|"RT @NotJoshEarnest: Listen up folks! Just because we lie about everything, doesn't mean we're lying about Russia hacking the election."
lovemrpibb2|rwindrem|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
lovemrpibb2|nbcnews|0.0772|0.128|0.731|0.142|RT @rwindrem: US intelligence community distressed at Trump's remarks re Russian hack of US election.  Our story. https://t.co/cpyE5AL7d6
ShammaBoyarin|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Iceis_|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
DuckmanMarla|HuffPostPol|0.0|0.0|1.0|0.0|"Donald Trump says it is ""ridiculous"" to say Russia intervened in the election on his behalf. https://t.co/JllElNGXI9 via @HuffPostPol"
DuckmanMarla|huffingtonpost|0.0|0.0|1.0|0.0|"Donald Trump says it is ""ridiculous"" to say Russia intervened in the election on his behalf. https://t.co/JllElNGXI9 via @HuffPostPol"
MikayesFiona|twitter|0.3612|0.0|0.898|0.102|Maybe next you &amp; McCain will be asking for election Do-Over like ex-CIA nut job Bob Baer. U ppl little too close to https://t.co/psK2pVnzNC
Cathy789|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
DailyAdams|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
raycholebunny|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
raycholebunny|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
JoeBeOne|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
JoeBeOne|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
shadavigm|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
xo_rosalee|Amberlynnjane15|-0.0279|0.17|0.664|0.166|"RT @Amberlynnjane15: If you decide to say we're not friends over who I supported in the election, then you clearly never respected me as yo"
ford_russell|andieiamwhoiam|0.5267|0.065|0.75|0.185|"RT @andieiamwhoiam: Sorry Lefties, Russians, recounts, aliens (the extraterrestrial kind)...you will never get a new election.  Trump won."
timothyworkman9|BreitbartNews|-0.822|0.434|0.495|0.071|RT @BreitbartNews: Why do Democrats want a war with Russia so badly? https://t.co/KfMP9vzZsu
timothyworkman9|breitbart|-0.822|0.434|0.495|0.071|RT @BreitbartNews: Why do Democrats want a war with Russia so badly? https://t.co/KfMP9vzZsu
AlexFedora|michaelianblack|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
AlexFedora|twitter|-0.3167|0.223|0.777|0.0|RT @michaelianblack: This. Whole. Election. Fucking. Stinks. Baaaaaaaaad. https://t.co/iUWejHTqL4
TwardowskiAK|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
TwardowskiAK|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
larsbaek|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
tmcmill81|Find_Me_Value|0.4404|0.0|0.734|0.266|RT @Find_Me_Value: Moffett: Towers attractive still (12-09-16) https://t.co/NQkqxxWXQM https://t.co/tHghdIJQ8T
tmcmill81|fiercewireless|0.4404|0.0|0.734|0.266|RT @Find_Me_Value: Moffett: Towers attractive still (12-09-16) https://t.co/NQkqxxWXQM https://t.co/tHghdIJQ8T
LOLatSJWs|hautedamn|-0.3384|0.252|0.63|0.118|@hautedamn also the same people that laughed at and mocked anyone suggesting the DNC could rig the election...aka fucking morons.
CNNfakenews|mtracey|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
CNNfakenews|cnn|-0.128|0.073|0.927|0.0|"RT @mtracey: Former CIA spooks running to CNN to demand ""a new election"" ... nothing to see here, folks https://t.co/JvUMybjpq8"
Ivana11117|Love_The_Donald|0.34|0.0|0.844|0.156|RT @Love_The_Donald: Homeland Security tied to attempted hack of Georgia's election database: Report https://t.co/y6csoEblbJ
Ivana11117|cnbc|0.34|0.0|0.844|0.156|RT @Love_The_Donald: Homeland Security tied to attempted hack of Georgia's election database: Report https://t.co/y6csoEblbJ
DistanceRun|DistanceRun|-0.4588|0.136|0.864|0.0|RT @DistanceRun: @aravosis @DavidCornDC Investigate the Orwellian data mining Co Trump used to cheat on the election Cambridge Analytica CA
UncommonTart|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Andyrguapo|DrJillStein|-0.3612|0.128|0.872|0.0|"RT @DrJillStein: Michigan's election is a ""hot mess"" because of antiquated state laws and a sloppy voting system. #RecountMI https://t.co/W"
Andyrguapo|t|-0.3612|0.128|0.872|0.0|"RT @DrJillStein: Michigan's election is a ""hot mess"" because of antiquated state laws and a sloppy voting system. #RecountMI https://t.co/W"
ErengwaM|zoomzoom130|0.0|0.0|1.0|0.0|RT @zoomzoom130: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean. https://t.co/zfWOq
ErengwaM|t|0.0|0.0|1.0|0.0|RT @zoomzoom130: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean. https://t.co/zfWOq
conservativelez|warnerthuston|-0.5647|0.173|0.753|0.073|"RT @warnerthuston: Liberals now say Russia was good enough to hack 50 states' election systems, but too stupid to hack a single Secretary o"
DTritsch|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
mamalocaz|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
KimbaGross|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
JoshGatewood|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
bldouglasjr|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
StevenNantz|PattyMurray|0.6124|0.0|0.737|0.263|"@PattyMurray Yes. Senator, please insist on a bipartisan investigation of Russian intervention in the 2016 presidential election."
burredea|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
widricbj197|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
llgwat|hiddenAmericans|0.3612|0.12|0.681|0.199|"RT @hiddenAmericans: Cavuto Rips Obama: Fox Didnt Win An Election, You Lost It#TrumpFirsts https://t.co/eGYXFvqdRG https://t.co/q0h90jK1qJ"
llgwat|hiddenamericans|0.3612|0.12|0.681|0.199|"RT @hiddenAmericans: Cavuto Rips Obama: Fox Didnt Win An Election, You Lost It#TrumpFirsts https://t.co/eGYXFvqdRG https://t.co/q0h90jK1qJ"
keanleathers|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
lionheart_erin|petitions|0.6523|0.0|0.764|0.236|PETION TO THE SUPREME COURT: Invalidate Election Results Of 2016-Order A New Election #NotMyPresident #TheResistance https://t.co/YkN0w1Dkrg
Judigal|RealEdMosca|-0.6705|0.234|0.766|0.0|RT @RealEdMosca: Obvious Russian hacking forced #CrookedHillary to ignore working class voters &amp; cost her electionCouldn't be her own arro
itsweezie|neilpX|-0.5423|0.17|0.83|0.0|"RT @neilpX: If McCain and Graham are able to expose the treason promulgated in the election, they will deserve to be heralded as American h"
bamilekeeavon|ZaynDiamonds|-0.4215|0.203|0.797|0.0|RT @ZaynDiamonds: 59% of their machines randomly broke on election day?  https://t.co/Xl0lmZ3BkH
bamilekeeavon|twitter|-0.4215|0.203|0.797|0.0|RT @ZaynDiamonds: 59% of their machines randomly broke on election day?  https://t.co/Xl0lmZ3BkH
sasyecat|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
sasyecat|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
yolisnampa|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
deb0815|nytopinion|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
deb0815|nytimes|-0.2732|0.116|0.884|0.0|RT @nytopinion: In Mr. Trump the Russians likely saw a stunningly ignorant and malleable political novice. https://t.co/0Zof9Cl4bT https://
JimFliesHigh|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
seenorseems|DougHenwood|0.296|0.0|0.804|0.196|RT @DougHenwood: Its ok to manipulate some elections https://t.co/h4ZNsWx1nU https://t.co/HeuenVGwVZ
seenorseems|observer|0.296|0.0|0.804|0.196|RT @DougHenwood: Its ok to manipulate some elections https://t.co/h4ZNsWx1nU https://t.co/HeuenVGwVZ
CheckingTheMath|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
CheckingTheMath|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
Bellalindafox|penultimatepen|0.4019|0.0|0.876|0.124|RT @penultimatepen: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co
Bellalindafox|t|0.4019|0.0|0.876|0.124|RT @penultimatepen: Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump via @politicususa https://t.co
shyaesthetic|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
shyaesthetic|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
fredricgstewart|Newsmax_Media|-0.6705|0.314|0.686|0.0|"Spicer: 'Zero' Proof Russia Tilted Election, Denies RNC Was Hacked https://t.co/KDfdkYQdiD #Newsmax via @Newsmax_Media"
fredricgstewart|newsmax|-0.6705|0.314|0.686|0.0|"Spicer: 'Zero' Proof Russia Tilted Election, Denies RNC Was Hacked https://t.co/KDfdkYQdiD #Newsmax via @Newsmax_Media"
Shrekopher|twitter|0.0|0.0|1.0|0.0|Russia did not hack the USA to manipulate the election. https://t.co/hnTQBbEqIW
geewhizpat|drspl5|-0.1007|0.227|0.59|0.183|"RT @drspl5: Election needs to be nullified. 5 weeks yo stop it.Takes care if Tillerson, Bolton, etc. Stop being PC and fight! Yes, I'm angr"
DixieUte|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
rphawg3150|NPR|0.0|0.0|1.0|0.0|"RT @NPR: NPR has independently confirmed the CIA's new assessment, which concludes that ""Russia was trying to tip the election to Trump."" h"
Serpentine202|2crazy4books2|0.0|0.0|1.0|0.0|RT @2crazy4books2: @Serpentine202 The CIA has proof. GOP conspired to suppress. https://t.co/UriwbWI930
Serpentine202|petitions|0.0|0.0|1.0|0.0|RT @2crazy4books2: @Serpentine202 The CIA has proof. GOP conspired to suppress. https://t.co/UriwbWI930
Urdnot123|PrisonPlanet|-0.3453|0.139|0.861|0.0|RT @PrisonPlanet: Russia interfered in the election! (no evidence).LEFT FREAKS OUT.Saudi Arabia provably bankrolled Clinton's campaign.
snap1949|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
snap1949||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
PaddyTopp|RepublicanChick|-0.1779|0.082|0.918|0.0|"RT @RepublicanChick: Liberals are accusing Russia of influencing the election. At the same time, liberals enabled citizens of other countri"
yamatoejam|ProgressiveShay|-0.7579|0.338|0.597|0.065|RT @ProgressiveShay: @kierobar THIS is scary as shit. They want to discredit the election. omg.
BJenerik|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
LillyRobinsons|POTUS|-0.4019|0.162|0.838|0.0|@POTUS @JoeBiden @SenFeinstein  @OversightDems Why does election count if we know it was hacked? #NoConfidence
Modus_Operand_|MarkSimoneNY|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
Modus_Operand_|nytimes|0.6486|0.093|0.633|0.274|RT @MarkSimoneNY: FBI investigation concludes there's no evidence that Russia tried to help Trump win the election: https://t.co/VreXCA4NIs
HotNostrilsrFun|trumpwrongworld|-0.296|0.104|0.896|0.0|RT @trumpwrongworld: There is no evidence Russia interfered with election. Saudi Arabia funds Clinton and the media is silent. #FAKENEWS#
M5B1tch|FaceTheNation|0.7506|0.0|0.709|0.291|"RT @FaceTheNation: ""You can't make this issue partisan. It is too important. A fundamental part of a democracy is a free and fair election."
JackDavisAZ|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
tleydn|mcuban|0.0|0.0|1.0|0.0|"@mcuban our ""first round draft pick"" not concerned that CIA asserts that Russia interfered with the US election. How is that not mortifying?"
YngHandsomeMfka|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
carolinelv|Stevenwhirsch99|0.0|0.0|1.0|0.0|RT @Stevenwhirsch99: The same people that told us Benghazi was because of a YouTube video are now trying to tell us that #RussianHackers st
SRTCBass90|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
TheyBecameBirds|bellhooks|0.6249|0.0|0.718|0.282|RT @bellhooks: is to embrace our global unity and united global resistance. #election #bellhooks #Trump
TheBoliBic|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
kaygrivas49|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
HRCNJVolunteers|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
HRCNJVolunteers||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
portialaw|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ninuhdiaz|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
ninuhdiaz|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Margare86751378|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
25thcenturygirl|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
ToriGlass|ericgarland|0.0|0.0|1.0|0.0|RT @ericgarland: Do you tell America the day after the election that Russia spearfished all of our think tanks in brazen fashion?
MattMurph24|VABVOX|-0.7184|0.25|0.75|0.0|"RT @VABVOX: I can't be the only reporter who finds it odd after months of claiming election was rigged, @BernieSanders has no comment on Tr"
lbersch|Slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
lbersch|slate|-0.34|0.146|0.854|0.0|RT @Slate: Key senators: Reports of Russian election meddling should alarm every American: https://t.co/O3nv3P6ts3 https://t.co/zFD04tOQRM
haytalrin|KarenSkeens2|0.0|0.0|1.0|0.0|@KarenSkeens2 if #Trump goes then #Pence has to go also bc he benefited from the election interference just as Trump did. Can't separate him
Tarkan291|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
MosesRoss|emigre80|-0.3802|0.217|0.662|0.121|"RT @emigre80: Both Trump and Sanders were delighted to cry ""rigged election!"" when they ran against Clinton.Now that there's evidence? *C"
NoGunsNoGulag|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
NoGunsNoGulag|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
Tylertas|MysteryVFXSuper|-0.1139|0.109|0.891|0.0|RT @MysteryVFXSuper: Hey Donnie... How come you don't want an investigation into Russian influence on election? Don't you want to prove you
EdMahalick|Mediaite|0.3612|0.0|0.837|0.163|@Mediaite American interests were compromised. The election was just the venue. It's time for unity in defense of all Americans.
ad0rkay|danversohara|0.0|0.0|1.0|0.0|RT @danversohara: Everyone around me: the election is over get over itMe: https://t.co/ykfoZyr5k2
ad0rkay|twitter|0.0|0.0|1.0|0.0|RT @danversohara: Everyone around me: the election is over get over itMe: https://t.co/ykfoZyr5k2
henryrodgersdc|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
henryrodgersdc|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
mattiOgreen|NateSilver538|0.5584|0.0|0.82|0.18|RT @NateSilver538: I'll put it like this: Clinton would almost certainly be President-elect if the election had been held on Oct. 27 (day b
evapaterson|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
Lesmitch529|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
sean_mp3|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
sean_mp3|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
Judah_Embassy|FRANCE24|-0.2263|0.221|0.621|0.159|"Gambian president rejects election results, demands fresh polls https://t.co/kUtHDpHPOn via @FRANCE24"
Judah_Embassy|france24|-0.2263|0.221|0.621|0.159|"Gambian president rejects election results, demands fresh polls https://t.co/kUtHDpHPOn via @FRANCE24"
WendyMarcinkie1|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
denise68wn|stevesilberman|-0.5423|0.149|0.851|0.0|"RT @stevesilberman: .@EricGarland's panoramic history of the Bad Mojo that resulted in the ""election"" of Trump. Tweetstorm for the ages. ht"
vonliesse|DaysOfTrump|0.0|0.0|1.0|0.0|RT @DaysOfTrump: Former UK Ambassador to Uzbekistan: I've met the person. It wasn't a Russian. It was an insider leaking the emails. https:
CrockerDon|stevesilberman|-0.5423|0.149|0.851|0.0|"RT @stevesilberman: .@EricGarland's panoramic history of the Bad Mojo that resulted in the ""election"" of Trump. Tweetstorm for the ages. ht"
ThuglyNast|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
Drez1723|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
ToriGlass|ericgarland|-0.296|0.099|0.901|0.0|RT @ericgarland: Do you come out the day after this totally weird-smelling abomination of an election with all its technical difficulties?
fall_sapphire|carlbernstein|-0.836|0.357|0.643|0.0|No. @carlbernstein tried to  ring the warning bell on each tv appearance BEFORE the election. Ratings whore cablene https://t.co/gEGmAvWjyV
fall_sapphire|twitter|-0.836|0.357|0.643|0.0|No. @carlbernstein tried to  ring the warning bell on each tv appearance BEFORE the election. Ratings whore cablene https://t.co/gEGmAvWjyV
GeorgeShanko|Snowden|0.0|0.0|1.0|0.0|"RT @Snowden: .@NYTimes once sat on facts that could change the 2004 election result, citing ""fairness."" Now CIA/FBI do the same. https://t."
GeorgeShanko||0.0|0.0|1.0|0.0|"RT @Snowden: .@NYTimes once sat on facts that could change the 2004 election result, citing ""fairness."" Now CIA/FBI do the same. https://t."
xseane|giffmacshane|0.3182|0.0|0.874|0.126|RT @giffmacshane: #ElectionFraud #RussiaHacking Please sign the petitionCall for a new election in wake of Russia's involvement https://t
xseane||0.3182|0.0|0.874|0.126|RT @giffmacshane: #ElectionFraud #RussiaHacking Please sign the petitionCall for a new election in wake of Russia's involvement https://t
Dezdrew|LindseyGrahamSC|0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
Dezdrew||0.0|0.0|1.0|0.0|"RT @LindseyGrahamSC: Joint statement with Senators McCain, Schumer, and Reed on reports Russia interfered with the 2016 Election. https://t"
cpizer|paulkrugman|0.296|0.0|0.694|0.306|RT @paulkrugman: Yep. Tainted election. https://t.co/PtimIiiy6x
cpizer|twitter|0.296|0.0|0.694|0.306|RT @paulkrugman: Yep. Tainted election. https://t.co/PtimIiiy6x
frozenmn|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
freeloosedirt|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
modernactivism|ABC|0.6369|0.0|0.704|0.296|@ABC The world's best cyber army doesnt belong to Russia https://t.co/WkYXk0gJVI
modernactivism|reuters|0.6369|0.0|0.704|0.296|@ABC The world's best cyber army doesnt belong to Russia https://t.co/WkYXk0gJVI
lavndrblue|linkis|0.0|0.0|1.0|0.0|https://t.co/q5uduX7pOi
OBrien41216022|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
mia_candace|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
martyrabkin|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
martyrabkin|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
edmik95|nytimesworld|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
edmik95|nytimes|0.1872|0.083|0.803|0.114|"RT @nytimesworld: Did Russia hack the election to elect Trump? The C.I.A. says yes, the F.B.I. is not sure. https://t.co/U3Q6Oe8Qfg https:/"
vonHerff|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
vonHerff|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
GeorgetteMcClel|Khanoisseur|0.296|0.0|0.856|0.144|RT @Khanoisseur: Since election top 5 banks added an eye-watering $200B in market capBank stocks highest since 12/2007 as they await Trum
conniebyr|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
conniebyr|change|0.0|0.0|1.0|0.0|RT @starfirst: President Obama: Time to Call for a New General Election! - Sign the Petition! https://t.co/pQJTN9QGm4 via @Change
rachaelji|freddiedeboer|0.34|0.0|0.888|0.112|"RT @freddiedeboer: The most striking, consistent aspect of post-election behavior from Democrats is the absolute refusal to engage in real"
critz_ccritz|petitions|0.0|0.0|1.0|0.0|SCOTUS: Invalidate Election Results Of 2016 - Order A New Election https://t.co/HeA7hI5RWP
cosmoksmom|ChicagoMGD|0.4767|0.0|0.853|0.147|RT @ChicagoMGD: @aliasvaughn @ezlusztig Reminder it isn't just the @CIA 16 other intelligence agencies had evidence of Russia's interferenc
llsmith2449|CRMunoz|-0.7983|0.393|0.607|0.0|@CRMunoz: Where's the outrage over the Russia hack? (opinion) - https://t.co/e8AT07y68K https://t.co/oLPmNDo4Q3 FAKE NEWS
llsmith2449|CNN|-0.7983|0.393|0.607|0.0|@CRMunoz: Where's the outrage over the Russia hack? (opinion) - https://t.co/e8AT07y68K https://t.co/oLPmNDo4Q3 FAKE NEWS
kostopoulos_d|ChicagoMGD|0.4767|0.0|0.853|0.147|RT @ChicagoMGD: @aliasvaughn @ezlusztig Reminder it isn't just the @CIA 16 other intelligence agencies had evidence of Russia's interferenc
JenniferLMeyer|kjacobsedits|0.4574|0.0|0.85|0.15|RT @kjacobsedits: Looking for a pro-women organization you can support in the wake of the election? Try @girlswritenow! https://t.co/YyljR7
JenniferLMeyer|t|0.4574|0.0|0.85|0.15|RT @kjacobsedits: Looking for a pro-women organization you can support in the wake of the election? Try @girlswritenow! https://t.co/YyljR7
solutionary52|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
solutionary52|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
janelleholmes20|DailyNewsBin|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
janelleholmes20|palmerreport|-0.4215|0.141|0.859|0.0|RT @DailyNewsBin: Jim Crow in Michigan: 87 vote machines broke in Americas blackest city on Election Day https://t.co/RSMGUS5BCq
StefanHayden|funder|0.0|0.0|1.0|0.0|RT @funder: Ex Agent: If CIA proves Russian interference-US should hold new elections #TrumpLeaks #RussianHackers #msnbc #amjoy https://t.c
StefanHayden||0.0|0.0|1.0|0.0|RT @funder: Ex Agent: If CIA proves Russian interference-US should hold new elections #TrumpLeaks #RussianHackers #msnbc #amjoy https://t.c
TerriLSelby|NotJoshEarnest|-0.2144|0.078|0.922|0.0|"RT @NotJoshEarnest: The proof is overwhelming that Russia hacked our election, but you'll just have to take our word for it because we're n"
hickorycreekof2|MagicRoyalty|0.2942|0.0|0.905|0.095|"RT @MagicRoyalty: On election night, Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! http"
GARYHARTMAN|armed-services|0.0|0.0|1.0|0.0|https://t.co/NMmXqaVkHD... https://t.co/Ty26XXzqAO
mainemama48|thehill|0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
mainemama48||0.675|0.0|0.716|0.284|"RT @thehill: Nate Silver: Clinton ""almost certainly"" would've won if election were before Comey's letterhttps://t.co/yTZdnv1uW3 https://t."
BloopJustSayin|AndyRichter|-0.0258|0.191|0.622|0.187|"RT @AndyRichter: Never forget that when shown substantial evidence that Russia hacked US election, @SenateMajLdr chose party over country."
larryglatt1|WalshFreedom|0.6662|0.085|0.672|0.243|RT @WalshFreedom: So wait...the CIA says Russia messed with our election to help Trump win and Trump attacks...the CIA?Not Russia? He goe
joannanoon|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
DanceMyVoice|Lee_in_Iowa|-0.1857|0.139|0.749|0.112|"RT @Lee_in_Iowa: @TheDemocrats We are a whole lot more interested in what you're going to do about the HACKED ELECTION! Grow a spine, dammi"
KatH_NY|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
leehlawrence|nytopinion|0.0|0.0|1.0|0.0|RT @nytopinion: Why would President-elect Trump object to a thorough bipartisan probe into Russian meddling? https://t.co/zDopY4Hcs0 https:
leehlawrence|nytimes|0.0|0.0|1.0|0.0|RT @nytopinion: Why would President-elect Trump object to a thorough bipartisan probe into Russian meddling? https://t.co/zDopY4Hcs0 https:
Gary_Davis_7807|usacsmret|-0.6119|0.192|0.808|0.0|RT @usacsmret: Obama claims our intel community totally missed the rise of ISIS but they are 100% correct in claiming the Russians rigged o
prairielive|SolidBlue2012|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
prairielive|t|0.2023|0.0|0.904|0.096|RT @SolidBlue2012: Trump faces first significant post-election pushback from Republicans over CIA report on Russia - LA Times https://t.co/
50linesonly|tteegar|-0.5242|0.232|0.67|0.098|RT @tteegar: BREAKING #RussianHackers made Hillary screech like an old crabby grandma &amp; lose the election!Nobody should be fooled! #Fak
Honey604|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
ivey__angel|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
ivey__angel|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
lmegordon|DavidYankovich|-0.296|0.109|0.891|0.0|RT @DavidYankovich: There is no Democrat/Republican side to the Russian influence in this election.You are either a patriot or a traitor.
Morosoph|kurteichenwald|0.2263|0.102|0.764|0.135|"RT @kurteichenwald: Fact: When it was announced that Trump had won the election, the Duma (lower house of Russian parliament) broke out in"
Eviljohna|MtnMD|0.0|0.0|1.0|0.0|"RT @MtnMD: RT @eileendefreest: #ImStillNotOver fact that Trump, Comey, and GOP Congress aren't in jail yet for allowing Russia to decide th"
donjuanw|cfahooligan|0.2023|0.067|0.833|0.099|RT @cfahooligan: @mtracey Have you seen it yet? Clintonite Trolls like @VABVOX are now accusing Sanders of being apart of the Russians rigg
haleybesser|birbigs|-0.0387|0.05|0.95|0.0|RT @birbigs: There's evidence that Russia swayed the U.S. election &amp; we're supposed to NOT talk about it constantly? I'm sorry but that's u
Bacalovx|Yascha_Mounk|-0.4019|0.119|0.881|0.0|"RT @Yascha_Mounk: German officials: Russia hacked Bundestag, released secret docs, will likely try to influence '17 election as in USA http"
itsweezie|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
ThatPersonEddie|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
ThatPersonEddie|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
mpostles|CmmnSnse1|0.4926|0.073|0.731|0.196|RT @CmmnSnse1: Please lets NOT forget Obama encouraged Illegals/foreigners to vote N this last election! How is that not an act of #Treason
markusg82|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
ThirtyMinuteAbs|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
oldmanbraun|WalshFreedom|0.7992|0.058|0.677|0.266|"RT @WalshFreedom: There's evidence Russia messed around with our election, but cuz our guy won, people on my side are ok with that?That's"
gasper_peg|TrumpsNewsDaily|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
gasper_peg|yahoo|0.0|0.0|1.0|0.0|RT @TrumpsNewsDaily: Trump on Russia meddling in US election: 'I don't believe it' https://t.co/Vvj0P3QTGw via @YahooNews
NVPeople|ndtv|0.0|0.0|1.0|0.0|Donald Trump On Russia Meddling In US Election: 'I Don't Believe It' https://t.co/NdoLV0FcW8 ^NDTV https://t.co/06094ydYU3
kenbod|GavinNewsom|0.4767|0.0|0.853|0.147|RT @GavinNewsom: Trump put down U.S. intelligence agencies rather than acknowledge Russia's involvement in the election. His priorities her
lackland50|CoryBooker|0.4588|0.0|0.81|0.19|RT @CoryBooker: I join urgent call for Congress to form bipartisan select committee to investigate Russian interference in election: https:
jonvankin|PinotYouDidnt|0.0|0.0|1.0|0.0|"RT @PinotYouDidnt: ""Why isn't Bernie talking publicly about Russian election interference?"" Really? C'mon, you know why: He benefited from"
_ThePage|ndtv|0.0|0.0|1.0|0.0|Donald Trump On Russia Meddling In US Election: 'I Don't Believe It' https://t.co/Q8hJwPDiRB ^NDTV https://t.co/58uiGO34DT
blueskymountain|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
rohitsh020678|Dev_Fadnavis|0.0|0.0|1.0|0.0|"RT @Dev_Fadnavis: Addressed today's first election campaign rally with @raosahebdanve ji at Gangapur in Aurangabad district, earlier today."
_dpaj|ndtv|0.0|0.0|1.0|0.0|Donald Trump On Russia Meddling In US Election: 'I Don't Believe It' https://t.co/oCjk9Q9lS0 ^NDTV https://t.co/ZJ3xB1hXEr
Emme69mw|cerenomri|0.0|0.0|1.0|0.0|"RT @cerenomri: Remember that one week during the election when the left was really, really concerned about anti-Semitism?They're supporti"
sunlightwarden|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
stksans|ABC|0.0|0.0|1.0|0.0|RT @ABC: NEW: Bipartisan group of senators release joint statement calling for examination of reports of Russian interference in 2016 US el
stanrails_store|twitter|0.0|0.0|1.0|0.0|Trump dismisses allegations of Russian election tampering; senators plan investigation - U.S. - Stripes https://t.co/1TpV6D4qPc
hailhail97|Steven_Strauss|-0.128|0.067|0.933|0.0|RT @Steven_Strauss: Trump: Obama is a Kenyan MuslimFox: America needs to hear this CIA: Putin tried to rig election for Trump Fox: we c
dcpatti13|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
Canada4TrumpNow|MarkSimoneNY|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
Canada4TrumpNow|twitter|-0.3612|0.2|0.8|0.0|RT @MarkSimoneNY: A picture of the people who rigged the election: https://t.co/Ma08WgVLko
TxsleuthUSA|cerenomri|0.0|0.0|1.0|0.0|@cerenomri Trump might not be POTUS if that had happened before election.
LanthaQ|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
LanthaQ|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
MahGill|morningmoneyben|-0.2263|0.112|0.888|0.0|@morningmoneyben I wonder if all of those Russian Twitter bots that disappeared after the election will return...
PSBbazmalea|YouTube|0.0|0.0|1.0|0.0|HAITI NEWS ELECTION 2016 TANDE KI SA Liliane Pierre Paul DI SOU ELECTION: https://t.co/OSCkwfDJuN via @YouTube
PSBbazmalea|youtube|0.0|0.0|1.0|0.0|HAITI NEWS ELECTION 2016 TANDE KI SA Liliane Pierre Paul DI SOU ELECTION: https://t.co/OSCkwfDJuN via @YouTube
M5B1tch|mhmck|0.0|0.0|1.0|0.0|"RT @mhmck: Rerun the election. Paper ballots. Two names: Clinton, Trump. International observers by the tens of thousands. Ukraine did it."
Marypat714|davebernstein|-0.4019|0.114|0.886|0.0|RT @davebernstein: Former CIA agent Robert Baer said any other country would hold a new election they found out they were hacked. (6/10)htt
SOcean5|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
RobbieGramer|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
ElizbethLManess|LeahR77|0.1531|0.11|0.758|0.133|RT @LeahR77: Lets Talk Foreign Govts Influencing An Election &amp; Bonus Getting Uranium &amp; Weapons Deals From SOS HRC For #FakeNews #Russians
DannyLinhardt|ParkerMolloy|-0.5067|0.17|0.83|0.0|"RT @ParkerMolloy: ""patrioteagle.flag says there's a child sex pizza dungeon!""""On it!""""The CIA says Russia messed w/ the election!""Some s"
ProvaxShill|AlyssaColeLit|-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
ProvaxShill||-0.4767|0.129|0.871|0.0|"RT @AlyssaColeLit: ""state officials are now admitting that most of the voting machines in Detroit were broken on Election Day"" Hmm. https:/"
anobscureartist|davebernstein|-0.4019|0.114|0.886|0.0|RT @davebernstein: Former CIA agent Robert Baer said any other country would hold a new election they found out they were hacked. (6/10)htt
2020pleasehurry|FaceTheNation|-0.0516|0.112|0.784|0.104|"RT @FaceTheNation: ""Russia tried to turn the election ... It means that Russia attacked the United States."" @TIME's Michael Duffy on CIA in"
foodnpolitics|businessinsider|0.5719|0.0|0.844|0.156|This article is a perfect example of why we've felt as if Earth has swung off its axis since Election Day: https://t.co/QVf8m7DCFs
ARayRobinson|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
SarahsMimi|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
SarahsMimi||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
Anyshka|GoddessKerriLyn|0.0|0.0|1.0|0.0|RT @GoddessKerriLyn: Rep. John Lewis submitted bill to Congress authorizing 2nd National ElectionPls call  your House reps 2 support!h
Chance32001459|Irwin_Elaine|0.0|0.0|1.0|0.0|RT @Irwin_Elaine: @_0HOUR1 Here's a list of all the Foreign Governments who interfered in the last Pres election. I mean... donated to the
billlm|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
beebecathy|MrJamesonNeat|-0.6597|0.231|0.769|0.0|RT @MrJamesonNeat: In states where election fraud seems rampant lawsuits should be filed to disqualify Trump electors @tribelaw @lessig htt
Jabulil20062214|jchaltiwanger|-0.0857|0.107|0.763|0.131|RT @jchaltiwanger: 60% of Americans supported Iraq invasion w/ NO EVIDENCE of WMDs. But NOW they want to see evidence to believe Russia int
KravSeattle|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
KravSeattle|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
SharonS72105601|trump_woman|0.0|0.0|1.0|0.0|RT @trump_woman: GOP Says CIA Must Show Evidence Russia Intervened In The Electionhttps://t.co/knQdr0iJC5 via @trump_woman #FakeNews #Jiha
SBace6|thehill|-0.34|0.217|0.616|0.167|"@thehill Is this the same @FBI that released the fake @HRC email scandal a week before the election? Yeah, they're certainly credible."
CyberRabid|KestrelArts|0.0|0.0|1.0|0.0|@KestrelArts @TrumpNewsUSA @6bird4 @CaroleDoms @nypost America goes 'red!' Proof that #RussiaHacking steered election.
HLNEditor|awakenedwire|0.0|0.0|1.0|0.0|Why the CIA Claims of Russian Interference in the U.S. Presidential Election Dont Make Sense https://t.co/zlGkeDLcba
JonRuhe|RogersParkMan|-0.3818|0.11|0.89|0.0|"RT @RogersParkMan: Hey @fakedansavage , think R's would be upset if Russians are found to have tampered with the R Primaries, not just the"
chloewweee|TopRopeTravis|0.6124|0.0|0.762|0.238|"RT @TopRopeTravis: Trump pre-election: We're going to #draintheswamp.Trump post-election: Just kidding, I'm hiring all of my rich buddies"
Fern0947|btstangel1|-0.1363|0.119|0.783|0.098|"@btstangel1 @Fern0947 @TIME @SugarMama7 Get over it, you LOST the election, move on, you're acting like a sour puss, a left wing nut bar."
kausikdatta22|stevesilberman|-0.5423|0.149|0.851|0.0|"RT @stevesilberman: .@EricGarland's panoramic history of the Bad Mojo that resulted in the ""election"" of Trump. Tweetstorm for the ages. ht"
CatholicGirl15|yahoo|0.0|0.0|1.0|0.0|"Nut! Trump slams 'ridiculous' report of Russian election hacking, claims Obama could be trying to unde... https://t.co/93hppMRQ1k via @yahoo"
CatholicGirl15|finance|0.0|0.0|1.0|0.0|"Nut! Trump slams 'ridiculous' report of Russian election hacking, claims Obama could be trying to unde... https://t.co/93hppMRQ1k via @yahoo"
AwakenedNews|awakenedwire|0.0|0.0|1.0|0.0|Why the CIA Claims of Russian Interference in the U.S. Presidential Election Dont Make Sense https://t.co/HBQ3B2QZwo
cardoc813|RanttNews|-0.34|0.146|0.854|0.0|RT @RanttNews: Russian interference in our election should alarm every American. We must dutifully reacthttps://t.co/FI0RjgEWmP
DLN_Editor|awakenedwire|0.0|0.0|1.0|0.0|Why the CIA Claims of Russian Interference in the U.S. Presidential Election Dont Make Sense https://t.co/CrxrOYixKd #durham
Goodnightma|RepublicanChick|-0.1779|0.082|0.918|0.0|"RT @RepublicanChick: Liberals are accusing Russia of influencing the election. At the same time, liberals enabled citizens of other countri"
stksans|twitter|-0.1531|0.063|0.938|0.0|"At this point, as more is revealed of his ties to Russia, the electors may have no choice but to call for new elect https://t.co/zAxzjtyzz0"
Maxbjaa|TheDailyEdge|-0.6597|0.293|0.579|0.128|"RT @TheDailyEdge: Trump tweets fake news from Infowars about election fraud, then puts Reince on TV to call CIA's best analysis an ""insane"
therussophile|therussophile|-0.4019|0.231|0.769|0.0|How To Instantly Tell If Russia Hacked theElection https://t.co/5i9WYA6Oyi https://t.co/XWIWhUhSoU
ASedlander|EJDionne|-0.5423|0.234|0.659|0.106|RT @EJDionne: Why a #Trump presidency inspires fear. My column: Russia's role in his election is scary. His response: Even more sohttps://
Bklyn2246|ezlusztig|0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
Bklyn2246||0.6124|0.103|0.676|0.221|RT @ezlusztig: That's it: FIVE. The rest of them are happy to have an enemy hack our democracy if it means they win an election. https://t.
J45553957J|alexanderhiggins|-0.6259|0.313|0.687|0.0|"This is what happened. An Attempt, but not successful https://t.co/AZ3Wzj3YfH"
Chande87|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
Sumenn7063|mattdpearce|-0.0516|0.096|0.816|0.089|RT @mattdpearce: Could you imagine the holy fit Trump would be throwing if there were signs China had hacked his staff to throw the electio
Hillary16IsBAE|ericgarland|0.0|0.0|1.0|0.0|RT @ericgarland: Do you tell America the day after the election that Russia spearfished all of our think tanks in brazen fashion?
TheeErin|markoff|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
TheeErin|t|-0.25|0.136|0.777|0.087|RT @markoff: Michigan officials admit majority of Detroit vote counting machines broke on Election Day - Palmer Report https://t.co/Gx9btLq
2crazy4books2|quinncy|-0.5093|0.397|0.603|0.0|@quinncy @BalmyBalmer @PalmerReport @DailyNewsBin Outrageous! https://t.co/UriwbWI930
2crazy4books2|petitions|-0.5093|0.397|0.603|0.0|@quinncy @BalmyBalmer @PalmerReport @DailyNewsBin Outrageous! https://t.co/UriwbWI930
natejgreen|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
weellio01|theguardian|0.5859|0.0|0.759|0.241|"FBI covered up Russian influence on Trump's election win, Harry Reid claims https://t.co/6j6g1iCN4c"
lopezpaul294|marcorubio|0.8074|0.0|0.7|0.3|RT @marcorubio: Congratulations to @JohnKennedyLA on winning his election today in Louisiana.  I look forward to our service together.  #LA
LivingNonActor|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
summerasana|VABVOX|0.0|0.0|1.0|0.0|"RT @VABVOX: .@SpeakerRyan is tweeting about overturning #Obamacare, not Russian interference with our election. https://t.co/4SirvxWCKi"
summerasana|twitter|0.0|0.0|1.0|0.0|"RT @VABVOX: .@SpeakerRyan is tweeting about overturning #Obamacare, not Russian interference with our election. https://t.co/4SirvxWCKi"
KathleenELoughr|DisavowTrump16|0.0|0.0|1.0|0.0|RT @DisavowTrump16: U.S. Concludes that Russia was involved in our election! RETWEET to to tell the Electoral College to vote for Hillary!
LikusPJ|JuddLegum|0.4404|0.0|0.847|0.153|RT @JuddLegum: Updated list of GOP members supporting investigation into Russian interference w/prez electionSen GrahamSen McCainSen Co
ActionTime|ActionTime|0.8455|0.0|0.663|0.337|RT @ActionTime: Please Retweet:All US Security Agencies Should FULLY Brief Every Member of Electoral College on How Russia Helped Trump WON
8802Ditman|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
greg_greer|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
YaoMingMtEverst|JohnWDean|0.0|0.0|1.0|0.0|RT @JohnWDean: The intel report on Russia's role in the 2016 election must be available for all electors before the electoral college meets
patriot_family|JBurtonXP|-0.4019|0.124|0.876|0.0|"RT @JBurtonXP: Always remember that by ""hacked the election,"" these people mean ""released 100% authentic documents that showed real Democra"
tzsawyer|JimGoldgeier|0.2732|0.0|0.909|0.091|"RT @JimGoldgeier: George HW Bush election in '88, the last time Democrats and Republicans alike accepted legitimacy of new POTUS, seems lik"
cathyboothfob|BreitbartNews|-0.1531|0.074|0.926|0.0|"RT @BreitbartNews: CORRECTION: After feedback from several Twitter folks, we now know there are NOT frequent food shortages in Ghana. https"
ZaynDiamonds|twitter|-0.4215|0.237|0.763|0.0|59% of their machines randomly broke on election day?  https://t.co/Xl0lmZ3BkH
dylanbailey7591|ericgarland|-0.4404|0.116|0.884|0.0|"RT @ericgarland: But from about 2009 to the 2016 election, a madness is being brewed and slowly poured down the throats of increasingly hys"
blueskymountain|blueskymountain|0.0|0.0|1.0|0.0|RT @blueskymountain: Ex-CIA operative calling for NEW Election: Any other country/democracy would.https://t.co/sCWpJ7stJD
lyndsay5SOS|KendallWellsx|0.8096|0.0|0.671|0.329|RT @KendallWellsx: I'm so ready to oust Wynne. Happy to be legally able to vote at the next Provincial election.
ClaireDiSalle|mashable|0.0|0.0|1.0|0.0|RT @mashable: The one social platform actually taking action ahead of Trump's America https://t.co/4Q3d2SnM5G https://t.co/41TlUUVzx2
ClaireDiSalle|mashable|0.0|0.0|1.0|0.0|RT @mashable: The one social platform actually taking action ahead of Trump's America https://t.co/4Q3d2SnM5G https://t.co/41TlUUVzx2
mackbarron|SarahPalinUSA|-0.0422|0.118|0.77|0.112|RT @SarahPalinUSA: Russia's getting out of hand? So says the defeated. Not to worry... remember I can keep an eye on them from here. https:
DMMadora|mitchellvii|-0.5574|0.195|0.805|0.0|RT @mitchellvii: So the Democrats are claiming that the Russians rigged the election by exposing what Democrats really think?You can't ma
mocheaptalk|Yascha_Mounk|-0.4019|0.119|0.881|0.0|"RT @Yascha_Mounk: German officials: Russia hacked Bundestag, released secret docs, will likely try to influence '17 election as in USA http"
magasouthern|TCB_AK|0.2942|0.0|0.905|0.095|RT @TCB_AK: On election night #Trump offered to buy Hillary's $7 million dollars worth of fireworks for 5 cents on the dollar! #Flashbac
kshark001|TimRunsHisMouth|0.0|0.0|1.0|0.0|RT @TimRunsHisMouth: Here's a list of all the Foreign Governments who interfered in the last Presidential election. I mean... donated to th
deejay90192|starfirst|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
deejay90192|msnbc|0.0|0.0|1.0|0.0|RT @starfirst: Wash Post: CIA concludes Russia interfered with 2016 election https://t.co/UpsdBNBRRk via @msnbc
NYpoet|TimOBrien|0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
NYpoet||0.296|0.109|0.698|0.194|"RT @TimOBrien: We're now in the era of a PEOTUS who dismisses facts, routinely lies, and creates false realities for supporters: https://t."
vicster|Shoq|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
vicster|t|0.4374|0.0|0.855|0.145|"RT @Shoq: THIS PETITION NEEDS 50 MILLION SIGNATURES, stat! Please pass it to everyone you've known since Kindergarten!https://t.co/XASXr"
takief|JuddLegum|0.4404|0.0|0.838|0.162|RT @JuddLegum: UPDATE: GOP members supporting investigation of Russian interference in electionSen GrahamSen McCainSen LankfordSen Cor
mortis_a|greenhousenyt|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
mortis_a|t|-0.25|0.151|0.753|0.097|RT @greenhousenyt: Michigan officials admit that a majority of Detroit's vote-counting machines broke on Election Day. https://t.co/GFLHaMg
TeresaMeyer2016|TheDemocrats|0.3612|0.0|0.894|0.106|RT @TheDemocrats: 2017 is going to be the most open and transparent DNC Chair election ever. Here's what that looks like: https://t.co/UuQm
TeresaMeyer2016|t|0.3612|0.0|0.894|0.106|RT @TheDemocrats: 2017 is going to be the most open and transparent DNC Chair election ever. Here's what that looks like: https://t.co/UuQm
2ALAW|steph93065|0.4215|0.0|0.887|0.113|"RT @steph93065: The same people that gave Hillary the debate questions &amp; got their ""news"" approved by Podesta are telling you Russia interf"
NancyOsborne180|tgreene319|0.5719|0.0|0.85|0.15|RT @tgreene319: Imagine if Clinton won amid intel that Russians interfered. GOP would have serial hearings &amp; Trump would Tweet hourly about
oufenix|MMFlint|0.8689|0.077|0.568|0.355|RT @MMFlint: The CIA has determined Russia hacked into our election to help elect Donald J. Trump. Now Trump names Putin best friend as OUR
ImDuchessK|thehill|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
ImDuchessK|twitter|0.0|0.0|1.0|0.0|RT @thehill: FBI breaks with CIA on Russian motives for interfering in U.S. electionhttps://t.co/iB3SfByyup https://t.co/byicz0v0lE
LEISUREGODDESS|JasonKander|-0.6597|0.213|0.787|0.0|"RT @JasonKander: If we ignore Russian espionage in our election, we embolden other foreign powers to launch similar attacks on every aspect"
DashieBotism|THEFATTESTCUNT|0.0|0.0|1.0|0.0|"@THEFATTESTCUNT This election was a sub, get me started on the fucking chavs."
dean_spagnoli|FitzyGFY|-0.7574|0.319|0.681|0.0|RT @FitzyGFY: I'm w/@mtdisme - Russia absolutely hacked into Steelers PSI last week to distract from US election accusations #DeflateGate2
LochTheScot|Miami4Trump|0.6833|0.14|0.594|0.266|"RT @Miami4Trump: Sorry Libs, Lindsey &amp; John Don't Qualify As Bilateral Support For Your BOGUS, Putin Hacked The Election Fairytale! LMAO "
Tankmanbrad|_Makada_|-0.8074|0.307|0.693|0.0|RT @_Makada_: The same fake news media who said it was impossible to rig the election are now claiming Russia rigged the election with no p
RedSoxNationMT|BreitbartNews|-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
RedSoxNationMT||-0.6124|0.306|0.603|0.091|"RT @BreitbartNews: 2016: When the ""pros"" accepted unconfirmed speculation as fact and demanded that politicians prove a negative. https://t"
anblanx|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
anblanx|washingtonpost|-0.3182|0.15|0.778|0.072|"RT @washingtonpost: Kellyanne Conway calls CIA report on Russian election meddling ""laughable and ridiculous"" https://t.co/SjxZTobti2"
irwin47shari|asamjulian|-0.34|0.193|0.714|0.092|"RT @asamjulian: Crazy Dem strategist suggests retaliation towards Russia for hacking our election, even though she admits theres no smok"
mariahorton14|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
mariahorton14|washingtonpost|-0.4588|0.235|0.765|0.0|"RT @washingtonpost: As Democrats demand probe over CIA election claim, GOP senators express doubt https://t.co/bWtLadv2Jm"
gilesgoatboy|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
monicalstone|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
LindsaySpell|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
blueskymountain|blueskymountain|0.7777|0.0|0.746|0.254|RT @blueskymountain: @drtommartinphd @52fairway Yes! So why is USA letting Russia win allowing trump to still be peotus?Why are we not rej
KellyLWilliams|SenJohnMcCain|-0.296|0.099|0.901|0.0|RT @SenJohnMcCain: #CyberSecurity can't be partisan. The stakes are too high. Will work across aisle to investigate &amp; stop cyberattacks htt
IqbalSharifBiru|twitter|0.4215|0.0|0.865|0.135|Donald J.Trump is The 45th Elect President of United States of America with a landslide victory.See my Facebook Act https://t.co/mAIRkrRa3h
mancari_brandy|Stevenwhirsch99|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
mancari_brandy|t|0.4005|0.0|0.876|0.124|RT @Stevenwhirsch99: Flashback to when Obama told Putin he would have more flexibility after the election. Catching on yet? https://t.co/xU
BillLonbeck|KellyannePolls|-0.3182|0.099|0.901|0.0|"RT @KellyannePolls: Now match the 1.2 billion dollars with the ""winning"" campaign messages and the post-election spin as to why they lost."
mgeneris|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: Another thing that isn't normal: there has not been a single moment since 11/8 where some part of me wasn't thinking a
Diortem|aston_wave|-0.4215|0.359|0.641|0.0|RT @aston_wave: I'm bitter: The Articlehttps://t.co/luqJotsJwS
DistractdMasses|BlackAutonomist|-0.5267|0.167|0.833|0.0|RT @BlackAutonomist: There is still no evidence of Russia rigging the US election. There is still no evidence of Russia rigging the US elec
damonbethea1|DavidYankovich|-0.296|0.109|0.891|0.0|RT @DavidYankovich: There is no Democrat/Republican side to the Russian influence in this election.You are either a patriot or a traitor.
naffis|pierre|0.5927|0.0|0.839|0.161|RT @pierre: Russia has Republican info but only released Democrats'. Can't imagine how holding on to it might be useful. https://t.co/SB4VX
naffis|t|0.5927|0.0|0.839|0.161|RT @pierre: Russia has Republican info but only released Democrats'. Can't imagine how holding on to it might be useful. https://t.co/SB4VX
SpacedSusan|michaelianblack|0.0|0.0|1.0|0.0|RT @michaelianblack: EITHER World's foremost intellgence agency is correct that Russia interfered in US election. ORDonald Trump is t
AriCostello|theguardian|-0.0258|0.196|0.613|0.19|Intelligence figures fear Trump reprisals over assessment of Russia election role https://t.co/iyYCc6SUht
SetthemF|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
PolarVan|Khanoisseur|0.0|0.0|1.0|0.0|"RT @Khanoisseur: Not only did Trump ask Russia to hack a political rival, he took millions from them before the election @1liners https://t"
PolarVan||0.0|0.0|1.0|0.0|"RT @Khanoisseur: Not only did Trump ask Russia to hack a political rival, he took millions from them before the election @1liners https://t"
hsummer|ChrisJZullo|0.0|0.0|1.0|0.0|"RT @ChrisJZullo: .@POTUS, still looking for post election plans? Run for a house seat with a 50 state ""Speaker of the House"" #flipthehouse"
hexogennotsugar|theonlyadult|-0.3164|0.098|0.902|0.0|RT @theonlyadult: The noise you just heard is the popping of a vein in my forehead. Cancel the fucking election results now! https://t.co/8
hexogennotsugar|twitter|-0.3164|0.098|0.902|0.0|RT @theonlyadult: The noise you just heard is the popping of a vein in my forehead. Cancel the fucking election results now! https://t.co/8
JeramySinopoli|ActionTime|0.6124|0.0|0.783|0.217|RT @ActionTime: Please Retweet:Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump #Resistance https:/
JeramySinopoli||0.6124|0.0|0.783|0.217|RT @ActionTime: Please Retweet:Calls Grow For A New Presidential Election To Be Held After Russia Meddled To Help Trump #Resistance https:/
xpro1|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
queene4theday|lpolgreen|0.7269|0.0|0.757|0.243|"RT @lpolgreen: I have covered many African elections. I have a pretty good idea how western election observers would respond to this in, sa"
lorilpeabody|KellyannePolls|0.0|0.0|1.0|0.0|"RT @KellyannePolls: FBI: ""fuzzy"", ""ambiguous"" connection. Did Putin's Russia really try and get Trump elected? CIA veterans urge caution ht"
ctpdenver|DavidYankovich|-0.296|0.109|0.891|0.0|RT @DavidYankovich: There is no Democrat/Republican side to the Russian influence in this election.You are either a patriot or a traitor.
dmendelsohnaviv|Steven_Strauss|-0.3612|0.194|0.711|0.095|"RT @Steven_Strauss: Man who thought HRC should lose security clearance over e-mail server, sees no need for investigation into Russian hack"
_zakaali|casatino|-0.1027|0.097|0.903|0.0|RT @casatino: FBI: sends vague letter; actually nothingMSM: *quivers*CIA: confirms Russia interfered w/electionMSM: \_()_/https://
