User|Original_User/Web|Compound|Negative|Neutral|Positive|Tweet
march4progress|Vallmeister|0.3182|0.0|0.892|0.108|RT @Vallmeister: Please take a moment to reflect on everything Bernie did for Equality and more Progressive policies during this election #
MacDHistory|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Police respond to shooting near Los Angeles-area polling place https://t.co/1255zj2WzQ
MacDHistory|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Police respond to shooting near Los Angeles-area polling place https://t.co/1255zj2WzQ
Dwtjr2|1VoiceMatters|-0.7793|0.327|0.673|0.0|RT @1VoiceMatters: This Election is RIGGED! This is unacceptable! #myvote2016 #ElectionDay #ElectionNight @bfraser747 @peddoc63 @_CFJ_ htt
glahn_|YouTube|0.0|0.0|1.0|0.0|Election Results and Analysis Live Stream https://t.co/LoBczIPoAv via @YouTube
glahn_|youtube|0.0|0.0|1.0|0.0|Election Results and Analysis Live Stream https://t.co/LoBczIPoAv via @YouTube
emily_jecker126|jolie_anderson9|0.5719|0.0|0.837|0.163|RT @jolie_anderson9: if Hilary wins the election she's gonna have to build a wall to keep us in bc I'm out
carlawinston5|Mrlend|0.5904|0.0|0.857|0.143|"RT @Mrlend: TELL ALL FRIENDS ESPEC FL, PA, VA, NC - GET OUT AND VOTE YOU'LL DECIDE ELECTION.. POLLERS SAY LATE VOTERS DECIDING = VOTE @TR h"
PattyHamilton19|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
silverfoxmedia1|kilmeade|0.7003|0.0|0.633|0.367|"RT @kilmeade: Special election edition of ""Kilmeade and Friends"" 7pm-9am https://t.co/gfZjqu8eBj  @foxandfriends"
silverfoxmedia1|radio|0.7003|0.0|0.633|0.367|"RT @kilmeade: Special election edition of ""Kilmeade and Friends"" 7pm-9am https://t.co/gfZjqu8eBj  @foxandfriends"
Sarklor|maragrunbaum|0.1406|0.0|0.925|0.075|"RT @maragrunbaum: Well, I came to the Botanical Garden this afternoon to try NOT to think about the election, but https://t.co/6ubdu4smf7"
Sarklor|twitter|0.1406|0.0|0.925|0.075|"RT @maragrunbaum: Well, I came to the Botanical Garden this afternoon to try NOT to think about the election, but https://t.co/6ubdu4smf7"
sillyri|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
wolfwood207|YouTube|0.4215|0.0|0.823|0.177|I liked a @YouTube video https://t.co/25urjYnm2g The Daily Show - The Final Days of the 2016 Election
wolfwood207|youtube|0.4215|0.0|0.823|0.177|I liked a @YouTube video https://t.co/25urjYnm2g The Daily Show - The Final Days of the 2016 Election
election_votes|C_Smatana|0.0|0.0|1.0|0.0|RT @C_Smatana: Who are you voting for Trump or Clinton?!? #ElectionDay #USElection2016 #ElectionNight #HillaryClintonForPresident #DonaldTr
mottstreet6|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
WHAS11NewsDesk|WHAS11Kayla|0.0|0.0|1.0|0.0|RT @WHAS11Kayla: Here's what KY Senate President Robert Stivers had to say ahead of tonight's election. The GOP has the... https://t.co/cCO
WHAS11NewsDesk|t|0.0|0.0|1.0|0.0|RT @WHAS11Kayla: Here's what KY Senate President Robert Stivers had to say ahead of tonight's election. The GOP has the... https://t.co/cCO
thatdaba|TheLastRefuge2|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
thatdaba|twitter|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
stratocat1012|Bikers4Trump|-0.6486|0.227|0.773|0.0|RT @Bikers4Trump: We need Trump &amp; #ImVotingBecause @HillaryClinton is a criminal &amp; must be stopped this Election Eve#RETWEET &amp; Visit https
BANQVE|Deggans|0.0|0.0|1.0|0.0|RT @Deggans: Follow #election 2016 results through NPR's live blog here: https://t.co/vcEZp5MQG1
BANQVE|npr|0.0|0.0|1.0|0.0|RT @Deggans: Follow #election 2016 results through NPR's live blog here: https://t.co/vcEZp5MQG1
awwhalenawl|iMustPandaLean|0.0|0.0|1.0|0.0|RT @iMustPandaLean: It's almost time for the results and I don't mean the election #CFP
SJB6991|bawesome84|0.9089|0.0|0.598|0.402|RT @bawesome84: Who do you honestly think will win the election? Not who you want to win but whom you think will win! @TinaCatalone @JtMobl
parettijacob|REALBrianStreng|0.7096|0.0|0.789|0.211|RT @REALBrianStreng: Joke is on Hillary if she wins the election because that means she has to sit at the desk Monica was under
EmmaSegasture|EpicallyKaren|-0.3472|0.238|0.617|0.144|RT @EpicallyKaren: #IVotedJillStein &amp; it felt so good to vote #PeoplePlanetAndPeaceOverProfit in this ridiculous insult of an election htt
JoeyVincent98|DrunkOldGrad|-0.481|0.135|0.865|0.0|RT @DrunkOldGrad: Here's a #MannequinChallenge from the Corps of Cadets to take your mind off this damn election for a minute. (Works cited
karodgers7|asuevents|0.6775|0.085|0.639|0.275|Check out this great event going on at ASU. Dont miss out! #Sponsored https://t.co/7AhPDQJYB1
tlynn561|kayleighmcenany|0.0|0.0|1.0|0.0|RT @kayleighmcenany: Evening voters could determine this election - you still have time to go vote Trump!!!  #ElectionNight
lilaustin110|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
blurrygambino|twitter|0.128|0.169|0.635|0.196|When you realize that we're screwed if trump or Hillary wins the election https://t.co/5ULRBFJVIR
RowenaGalavitz|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
RowenaGalavitz|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
M7MD_2oo1|IHE_OFFICIAL|-0.8625|0.312|0.688|0.0|"RT @IHE_OFFICIAL: I have a new video finished, but I'm thinking about saving it till all the election stress has died down a little."
mlynne3|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
sean_lynch|twitter|0.4019|0.0|0.891|0.109|"When Obama got elected, iPhone had been on sale for a year and had just added 3G support. Can't wait to see where c https://t.co/WMqj1zV2Ey"
freddie1012|Things4WhitePpl|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
freddie1012|twitter|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
SteveTVNews|secstatewa|0.0|0.0|1.0|0.0|RT @secstatewa: Here's how WA election returns will be reported tonight &amp; in coming days. https://t.co/BwDLwX4ING
SteveTVNews|twitter|0.0|0.0|1.0|0.0|RT @secstatewa: Here's how WA election returns will be reported tonight &amp; in coming days. https://t.co/BwDLwX4ING
See_My_Vest|fakedansavage|-0.2579|0.165|0.733|0.102|RT @fakedansavage: I'm retweeting a Republican without sarcasm or snark - this election is insane. https://t.co/mvaoZO0elr
See_My_Vest|twitter|-0.2579|0.165|0.733|0.102|RT @fakedansavage: I'm retweeting a Republican without sarcasm or snark - this election is insane. https://t.co/mvaoZO0elr
Zackdjohnson1|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
Zackdjohnson1|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
wolfwood207|YouTube|0.0|0.0|1.0|0.0|I added a video to a @YouTube playlist https://t.co/25urjYnm2g The Daily Show - The Final Days of the 2016 Election
wolfwood207|youtube|0.0|0.0|1.0|0.0|I added a video to a @YouTube playlist https://t.co/25urjYnm2g The Daily Show - The Final Days of the 2016 Election
aaronevaughn|ralphDrussoAP|0.0|0.0|1.0|0.0|"RT @ralphDrussoAP: Election Day. Or as sports writers call it, the day the news desk gets pizza for doing what the sports desk does every n"
nafi9918|SputnikInt|0.0|0.0|1.0|0.0|RT @SputnikInt: LIVE UPDATE: @realDonaldTrump currently leads @HillaryClinton as first polls close https://t.co/oTa25kErgX #USElection2016
nafi9918|sputniknews|0.0|0.0|1.0|0.0|RT @SputnikInt: LIVE UPDATE: @realDonaldTrump currently leads @HillaryClinton as first polls close https://t.co/oTa25kErgX #USElection2016
InfoOcheph|digitaltrends|0.3818|0.0|0.809|0.191|Electionland Google Trends map helps voters visualize polling station issues https://t.co/tNLOCfzT7D https://t.co/eY2c5VFy8E
SaltireComic|SaltireComics|-0.5178|0.143|0.857|0.0|RT @SaltireComics: Stressed out by Election Day? Need to know Scotland's got your back?Well we do! Check out our #ElectionDay deal!https:
Ali_leyva12|DanaiGurira|0.783|0.0|0.567|0.433|RT @DanaiGurira: Happy Election Day!Make sure your voice is heard!Vote!#ImWithHer.#TheFutureisFemale https://t.co/s6XK0ZYDzt
Ali_leyva12|twitter|0.783|0.0|0.567|0.433|RT @DanaiGurira: Happy Election Day!Make sure your voice is heard!Vote!#ImWithHer.#TheFutureisFemale https://t.co/s6XK0ZYDzt
CapeMayMeg|billy_penn|0.3412|0.0|0.862|0.138|RT @billy_penn: Some voting machines went down today. @Commish_Schmidt says don't worry about it. https://t.co/YDhwXcpWA6 https://t.co/CVcu
CapeMayMeg|billypenn|0.3412|0.0|0.862|0.138|RT @billy_penn: Some voting machines went down today. @Commish_Schmidt says don't worry about it. https://t.co/YDhwXcpWA6 https://t.co/CVcu
sethjpierce|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
ardie2pt0|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
ardie2pt0|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
LeighaCrumpler|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
LeighaCrumpler|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
CarpeMors90|JeniSelke1|0.4019|0.0|0.863|0.137|RT @JeniSelke1: @LeTHaLMiGRaiNe @JamesMArcher @SusanSarandon this is more than a single election. We are building a party for the people. #
Herityalia|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
Herityalia|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
sheacollagen|uniqueprophet|0.0258|0.153|0.691|0.157|"RT @uniqueprophet: OOPS @realDonaldTrump, @trump TRUMP SUPPORTERS, WE HAVE ENDURED TOO MUCH STRESS, EMOTION,EFFORT,DON'T LET LEFT SCUM STEA"
PacifierGaga|HuffingtonPost|0.0|0.0|1.0|0.0|RT @HuffingtonPost: 30 oddly insightful quotes from kids about the election https://t.co/0WwtoflHHU https://t.co/2ghyhcKAOh
PacifierGaga|m|0.0|0.0|1.0|0.0|RT @HuffingtonPost: 30 oddly insightful quotes from kids about the election https://t.co/0WwtoflHHU https://t.co/2ghyhcKAOh
Michael_Rokicki|yankeeclassic46|0.4404|0.0|0.854|0.146|"@yankeeclassic46 I wanted to watch Santos/Vinick election day episode to feel better. But, Leo. That would make it https://t.co/MErJPgCyXR"
Michael_Rokicki|twitter|0.4404|0.0|0.854|0.146|"@yankeeclassic46 I wanted to watch Santos/Vinick election day episode to feel better. But, Leo. That would make it https://t.co/MErJPgCyXR"
TwinParasite|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
TwinParasite|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
GrimKarl|LeahR77|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
GrimKarl|breitbart|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
stanleydob|twitter|0.6369|0.0|0.826|0.174|#FOXNEWS2016 Me and my pops watching the best election coverage on Fox News after both doing our part voting pro-li https://t.co/XSgV7HdHgo
agent_it|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
mayaventura_|twitter|0.0|0.0|1.0|0.0|"just goes to show you, this election isn't Democrats vs. Republicans. it's Those With Common Sense vs. Idiots https://t.co/m0iN450pwO"
FdeFossard|MujatiBrewing|-0.7096|0.396|0.604|0.0|Watching old vlogs by @MujatiBrewing to avoid all this election misery.
TRINITYPRAISE|mike_pence|0.0|0.0|1.0|0.0|"RT @mike_pence: This Election Day, America is standing at the crossroads of history. RT this if you're voting for @realDonaldTrump. Togethe"
outdoortechie|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
outdoortechie|t|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
CorianderSleuth|pardonbeggar|0.4404|0.0|0.854|0.146|RT @pardonbeggar: [doing standup]this election is truly neck and neckunfortunately one of the candidates is a giraffe::they take away
1blessedbee|healthandcents|-0.41|0.215|0.671|0.113|"RT @healthandcents: @payao1a1 ABSOLUTE TRUTH. If #Trump does not win this, we will never have free election again. #Globalists will control"
jodybufkin|MlquToast|0.7263|0.0|0.711|0.289|"RT @MlquToast: Election Night at #LimerickJunction Free comedy, drink deals, and the future of America! 10PM #atlcomedy"
DreamStarrCEO|MARLIT0|-0.0772|0.248|0.526|0.226|RT @MARLIT0: This election is an insult to intellect
TheHumpty|davidsirota|0.7351|0.0|0.828|0.172|"RT @davidsirota: I know Im going out on a limb here, but Im just gonna predict that the winner of the 2016 election will be money and cor"
dorriedeakins|DonaldJTrumpJr|0.3164|0.0|0.906|0.094|RT @DonaldJTrumpJr: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERSGET OUT AND VOTE! Find 5 others. This is our chance to take back Am
Cricaholics|itvnews|0.0|0.0|1.0|0.0|RT @itvnews: US Election: Stark difference between how men and women are expected to vote #Election2016 #ElectionNight https://t.co/BfQPcj2
Cricaholics|t|0.0|0.0|1.0|0.0|RT @itvnews: US Election: Stark difference between how men and women are expected to vote #Election2016 #ElectionNight https://t.co/BfQPcj2
janjeffcoat|instagram|0.0|0.0|1.0|0.0|Election Night... she just wants to watch #docmcstuffins &amp; Mommy has to go  for a 2 a.m. https://t.co/BMsWbJARCc
lyndacsmith|Stonewall_77|0.0|0.0|1.0|0.0|RT @Stonewall_77: BREAKING: Comey To Be Firedhttps://t.co/qq9ow5pCVQ#MAGA #TrumpTrain#ElectionDay https://t.co/7yRAvM78ba
lyndacsmith|twitter|0.0|0.0|1.0|0.0|RT @Stonewall_77: BREAKING: Comey To Be Firedhttps://t.co/qq9ow5pCVQ#MAGA #TrumpTrain#ElectionDay https://t.co/7yRAvM78ba
sgunn|ericasmith|0.0|0.0|1.0|0.0|RT @ericasmith: .@travislylesnews and @CatGRog are going to be snapping presidential election results tonight for @virginianpilot. Follow a
irisheyes8701|WDFx2EU8|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
irisheyes8701|t|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
BillWarp9|CNNPolitics|0.5719|0.0|0.802|0.198|"RT @CNNPolitics: BREAKING: Clinton wins traditional midnight vote in Dixville Notch, New Hampshire https://t.co/fVi0JzyFOr #CNNElection htt"
BillWarp9|cnn|0.5719|0.0|0.802|0.198|"RT @CNNPolitics: BREAKING: Clinton wins traditional midnight vote in Dixville Notch, New Hampshire https://t.co/fVi0JzyFOr #CNNElection htt"
LANDoCUH|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
LANDoCUH|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
Yad_FPEnergy|fpinvesting|0.1027|0.0|0.915|0.085|"Stocks, Canadian dollar and Mexican peso climb as investors await U.S. election results https://t.co/hD2b2owUo8 via @fpinvesting"
Yad_FPEnergy|business|0.1027|0.0|0.915|0.085|"Stocks, Canadian dollar and Mexican peso climb as investors await U.S. election results https://t.co/hD2b2owUo8 via @fpinvesting"
SAIS_MIEF|JHU_BIPR|0.0|0.0|1.0|0.0|"RT @JHU_BIPR: On #USElection2016, after @Erik_Jones_SAIS's introduction on the US Electoral College, a student panel discusses the effects"
bristyIes|G_Eazy|0.7644|0.0|0.752|0.248|"RT @G_Eazy: PLEASE GO OUT AND VOTE WHATEVER YOU DO, THIS COULD BE THE MOST IMPORTANT ELECTION OF OUR LIVES #imwithher #fuckdonaldtrump"
Darksbane7|SWatercolour|0.3182|0.0|0.881|0.119|RT @SWatercolour: My university is showing the election results at a student bar ending at 5am pray for me
paulwatermusic|jgillie302|0.0|0.0|1.0|0.0|RT @jgillie302: This election has been the EPITOME of House of Cards.#ElectionDay
StephenPoore804|YahooSports|0.0|0.0|1.0|0.0|RT @YahooSports: Ric Flair voted for exactly who you'd think Ric Flair would vote for: Ric Flair. https://t.co/2GceP31bit https://t.co/wI6G
StephenPoore804|sports|0.0|0.0|1.0|0.0|RT @YahooSports: Ric Flair voted for exactly who you'd think Ric Flair would vote for: Ric Flair. https://t.co/2GceP31bit https://t.co/wI6G
jimmybelshe|DRUDGE_REPORT|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
jimmybelshe|businessinsider|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
bear_oyo|ProfessorF|0.8225|0.0|0.703|0.297|"RT @ProfessorF: Wow another example of Hillary's ""superior"" ground game. That's brilliant. Having election officials tell people who to vot"
SMLongmate|BuzzfeedNews|0.6948|0.0|0.771|0.229|@BuzzfeedNews I am so happy you are reporting on the election  You guys are making this day bearable 
asahi_azumane|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
asahi_azumane|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
zaraki921|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
zaraki921|t|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
_LookDontTouch|blackvoices|0.5719|0.0|0.791|0.209|RT @blackvoices: Twitter turned election day into #ObamaDay to celebrate the first family https://t.co/vwUSM6Twom https://t.co/KpmapCx1pk
_LookDontTouch|huffingtonpost|0.5719|0.0|0.791|0.209|RT @blackvoices: Twitter turned election day into #ObamaDay to celebrate the first family https://t.co/vwUSM6Twom https://t.co/KpmapCx1pk
okayykaylaaa|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
CELEBUZZ|celebuzz|0.0|0.0|1.0|0.0|All of these celebrities voted. (Have you?) See a gallery of their voting selfies: https://t.co/ylspzRVx9c https://t.co/nvrkkiywcv
BestFrenz|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
BestFrenz|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
Sixkiller1835|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
twlldun|whoislukecusick|0.0|0.0|1.0|0.0|@whoislukecusick @youngvulgarian I sneakily unretweeted days ago to prepare for election night.
mushoe01|electionprojection|0.0|0.0|1.0|0.0|2016 Presidential election projections https://t.co/XsDzlPJXNu
Professor3535|TamEdwards6abc|0.4939|0.0|0.862|0.138|"RT @TamEdwards6abc: Women are flocking to Susan B Anthony's NY State gravesite, leaving their ""I Voted"" stickers on headstone, in honor of"
tennisballbondi|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
tennisballbondi|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
cbooooob|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
nemchocke|KellyScaletta|0.4019|0.0|0.856|0.144|"RT @KellyScaletta: ""Active shooter situation"" is NOT something we should see on election day. It's beyond despicable."
superjaberwocky|eidietrich|0.0|0.0|1.0|0.0|RT @eidietrich: Hot take from @TheOnion on Montana's role in the presidential contest. HT @CarterTroy https://t.co/r6qISw9lYx
superjaberwocky|theonion|0.0|0.0|1.0|0.0|RT @eidietrich: Hot take from @TheOnion on Montana's role in the presidential contest. HT @CarterTroy https://t.co/r6qISw9lYx
FM1888|Bro_Pair|0.0258|0.0|0.936|0.064|@Bro_Pair  I think my ceaseless tweeting about the election to my 140 porn-bot followers has prevented a Trump victory.
vancouverstuart|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
wvpe|npr|0.0|0.0|1.0|0.0|Explore online results while listening to 88.1 WVPE Public Radio https://t.co/wUtnOPMt4D
cdbarker|stefanielaine|0.8478|0.0|0.545|0.455|"@stefanielaine Hey, this is our first election night as like, friends, this is fun!"
Whyatt|CAC_ACE|0.7102|0.0|0.753|0.247|@CAC_ACE Making Ethical Decision @SoccerNS BMO Facility. Somewhat funny that this is being offered on the eve of th https://t.co/RhojWX4Oqr
Whyatt|twitter|0.7102|0.0|0.753|0.247|@CAC_ACE Making Ethical Decision @SoccerNS BMO Facility. Somewhat funny that this is being offered on the eve of th https://t.co/RhojWX4Oqr
NetflixChili|ComplexMag|0.0|0.0|1.0|0.0|RT @ComplexMag: We're live blogging the series finale of Americajoin us! https://t.co/UYu2z42U0g https://t.co/A2QXki1sar
NetflixChili|complex|0.0|0.0|1.0|0.0|RT @ComplexMag: We're live blogging the series finale of Americajoin us! https://t.co/UYu2z42U0g https://t.co/A2QXki1sar
markjonesaudio|ContenderGame|0.75|0.113|0.543|0.344|RT @ContenderGame: All domestic shipping at TheContender.us is FREE today! Treat yourself for surviving this insane election! Code: Election
FearDept|sexbsex|-0.5114|0.276|0.575|0.149|RT @sexbsex: Lmao people are so brainwashed they get so scared. What a fear induced election. Ah almost done....
tdoyle_86|MannieMforever|-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
tdoyle_86||-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
Amac_16|immigrant4trump|0.7506|0.0|0.766|0.234|"RT @immigrant4trump: If you make this go viral, Trump will win. It's about 2 minutes that makes the choice in this election crystal clear h"
PARGANEXTDOOR_|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
PARGANEXTDOOR_|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
JacobAClark13|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
JacobAClark13|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
FAOUOfficial|twitter|0.3612|0.0|0.667|0.333|Gary watching the election like https://t.co/De5EWO7hp8
lunaazul70|t|0.0|0.0|1.0|0.0|"https://t.co/64CmtER4LyLive coverage: Election Day 2016 coverage with Katie Couric, Matt Bai"
JebLadat|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
teokee|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: This election my dad did not spend time raising $ from the billionaire elite. Instead he spent time talking to the Amer
waterfunus43|DonaldJTrumpJr|-0.3595|0.098|0.902|0.0|RT @DonaldJTrumpJr: Media elites have done everything they can to stop Trump. WE THE PEOPLE will rise up and take back America! #Trump #Ele
Meganwiley204|DonaldJTrumpJr|-0.3595|0.098|0.902|0.0|RT @DonaldJTrumpJr: Media elites have done everything they can to stop Trump. WE THE PEOPLE will rise up and take back America! #Trump #Ele
von_non_|FareedZakaria|0.3612|0.0|0.783|0.217|@FareedZakaria would you like to get in an election prediction?
BrettSpielberg|netsirk12|0.3818|0.097|0.709|0.194|"RT @netsirk12: It's Election Day. Regardless of the outcome, I hope and pray that I never have to hear ""Fight Song"" ever again. #ElectionDay"
sofiafromkorea|rollcall|0.0|0.0|1.0|0.0|RT @rollcall: We're 2 hours away from the first set of major poll closings. How to watch election night: https://t.co/Bx1NZhAGPH https://t.
sofiafromkorea|rollcall|0.0|0.0|1.0|0.0|RT @rollcall: We're 2 hours away from the first set of major poll closings. How to watch election night: https://t.co/Bx1NZhAGPH https://t.
jjrbs|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
jjrbs|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
MaryEBarnes|goodtobeme0|0.0|0.0|1.0|0.0|RT @goodtobeme0: @goodtobeme0 States Poll Prediction of Election 2016 11/07/2016(Final)                  https://t.co/glH58Brt0W  @StatesPo
MaryEBarnes|twitter|0.0|0.0|1.0|0.0|RT @goodtobeme0: @goodtobeme0 States Poll Prediction of Election 2016 11/07/2016(Final)                  https://t.co/glH58Brt0W  @StatesPo
sueludad|HuffPostPol|0.4215|0.147|0.58|0.272|RT @HuffPostPol: This election was colossally dumb and we're all lucky we survived it https://t.co/xFLKuRqNmn https://t.co/OiHLgURoiC
sueludad|m|0.4215|0.147|0.58|0.272|RT @HuffPostPol: This election was colossally dumb and we're all lucky we survived it https://t.co/xFLKuRqNmn https://t.co/OiHLgURoiC
natsaysmiaow|carolineplz|-0.128|0.171|0.717|0.112|RT @carolineplz: Just got off the phone from a few Australian interviews-- weirdly comforted that they are also nervous about our election
melodicwaffle|stupeoscientia|0.0|0.0|1.0|0.0|RT @stupeoscientia: it's election day https://t.co/9HyCHL28xr
melodicwaffle|twitter|0.0|0.0|1.0|0.0|RT @stupeoscientia: it's election day https://t.co/9HyCHL28xr
twinkIouis|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
twinkIouis|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
mayadiez|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
abetrve|Suxting|0.3182|0.0|0.685|0.315|RT @Suxting: I've got a huge election.
andreww__14|MattMoretta|0.8934|0.0|0.545|0.455|"RT @MattMoretta: Plot twist: Matthew McConaughey wins election, everyone receives a brand new Lincoln, happiness is restored alright alrigh"
TeddyObo|Forbes|-0.6369|0.245|0.755|0.0|RT @Forbes: A nationwide election cyber attack is near impossiblebut these states are at risk of hacking: https://t.co/tiu0nhsMfa https://
TeddyObo|forbes|-0.6369|0.245|0.755|0.0|RT @Forbes: A nationwide election cyber attack is near impossiblebut these states are at risk of hacking: https://t.co/tiu0nhsMfa https://
Bassmavrik|JamesOKeefeIII|-0.4767|0.119|0.881|0.0|RT @JamesOKeefeIII: We'll have teams everywhere tomorrow. If you are doing something wrong on Election Day we find you we film you and we w
TheMadHessian|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
TheMadHessian|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
breaunaclifford|CALUMDATING|0.1571|0.115|0.737|0.147|RT @CALUMDATING: bless calum for tweeting about the election/voting even though he's not American + on holidays
JanayeMcGrew|JanayeMcGrew|0.814|0.0|0.624|0.376|@JanayeMcGrew what I'm saying is that I'd like to make Election Night fun and not scary again.
Kaori_2020|sugoibrooks|-0.1027|0.072|0.928|0.0|RT @sugoibrooks: Everyone's talking about the election while i'm getting shook over a 25 year old in a tigger onesie. https://t.co/IvsASgAJ
Kaori_2020|t|-0.1027|0.072|0.928|0.0|RT @sugoibrooks: Everyone's talking about the election while i'm getting shook over a 25 year old in a tigger onesie. https://t.co/IvsASgAJ
wiseguysliquors|instagram|0.5994|0.099|0.583|0.318|"No matter the outcome of this election, the Wise Guys crew encourages YOU to keep on https://t.co/VmhbLA7U7L"
MadAsis|SkyWilliams|0.0|0.0|1.0|0.0|RT @SkyWilliams: anyone got the Presidential Election Series Finale spoilers? 
KortKneee_Rae|twitter|0.0|0.0|1.0|0.0|It will serve as a much needed break from election results! I think it's going to be a longgggg night! #MarriedLife https://t.co/PIX0MRyh8T
HigashiNY|dril|0.0|0.0|1.0|0.0|RT @dril: if you ask me this election could end about 100 different ways:1) trump gets 0% of the vote2) trump gets 1% of the vote3) trum
JuliaaBlando|mallorywiest_|-0.128|0.16|0.71|0.13|RT @mallorywiest_: these arguments are almost as big of a joke as this election is
KatelynBruzzi|TheVoiceBHS|-0.4215|0.141|0.859|0.0|RT @TheVoiceBHS: Blackman High School's 2016 Mock Election Results for your comparison to the real election results https://t.co/DlMI2GPXMw
KatelynBruzzi|twitter|-0.4215|0.141|0.859|0.0|RT @TheVoiceBHS: Blackman High School's 2016 Mock Election Results for your comparison to the real election results https://t.co/DlMI2GPXMw
TheTruthhTeller|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
TheTruthhTeller|t|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
CloreenBacNSkin|dailydot|0.296|0.0|0.833|0.167|"RT @dailydot: Surviving 2016: Live election results, memes, and news: https://t.co/8Q2q2yU9LY https://t.co/CxX2Ml1bMc"
CloreenBacNSkin|dailydot|0.296|0.0|0.833|0.167|"RT @dailydot: Surviving 2016: Live election results, memes, and news: https://t.co/8Q2q2yU9LY https://t.co/CxX2Ml1bMc"
jeanne_tall|Caveman2743|0.4466|0.0|0.827|0.173|"RT @Caveman2743: RED ALERT: On Eve of Election, Benghazi BOMBSHELL Rains Down on Hillary https://t.co/rGox20vXgM"
jeanne_tall|conservativetribune|0.4466|0.0|0.827|0.173|"RT @Caveman2743: RED ALERT: On Eve of Election, Benghazi BOMBSHELL Rains Down on Hillary https://t.co/rGox20vXgM"
Witt_less00|livvylu582|0.7096|0.0|0.789|0.211|RT @livvylu582: This election will be like ripping off a bandaid but instead of relief you just realize that the wound didn't heal one bit.
oliviaisfake|carwash54|0.7085|0.0|0.734|0.266|"RT @carwash54: Me @ the beginning of the election: Ain't no way America letting a cheeto become president. lol what a joke Me November 7,"
CraftyOldFox|leighsales|0.0|0.0|1.0|0.0|RT @leighsales: Journos keep your eyes peeled for news that politicians and others try to bury after about 2pm this arvo as the US election
angelrains|video|0.4019|0.0|0.649|0.351|Donald Trump Election Watch Party | https://t.co/xvzumoMGWs
samanthrusso|twitter|0.4404|0.0|0.734|0.266|the only bright side to this entire election https://t.co/TThw8yoHxf
WavyKirk|FiveThirtyEight|0.4215|0.0|0.763|0.237|RT @FiveThirtyEight: Why Clinton is favored in Virginia. #ElectionNight https://t.co/QAF08CtpPW
WavyKirk|fivethirtyeight|0.4215|0.0|0.763|0.237|RT @FiveThirtyEight: Why Clinton is favored in Virginia. #ElectionNight https://t.co/QAF08CtpPW
shaycode|jason_howerton|-0.8481|0.365|0.635|0.0|"RT @jason_howerton: UPDATE: At least 1 dead, 3 injured in Azusa shooting, @latimes reports. Police dealing with heavily armed suspect: http"
biebrvogue|twitter|0.0|0.122|0.756|0.122|im actually tearing up bc this election is basically over and it's finally hitting me tht u didn't win ffs dammit t https://t.co/MIRPkGYGK4
meghiraki|carwash54|0.7085|0.0|0.734|0.266|"RT @carwash54: Me @ the beginning of the election: Ain't no way America letting a cheeto become president. lol what a joke Me November 7,"
mikaylacavenas|comedyandtruth|0.0|0.0|1.0|0.0|RT @comedyandtruth: Twitter on Election Day https://t.co/R3ihQKTfvr
mikaylacavenas|vine|0.0|0.0|1.0|0.0|RT @comedyandtruth: Twitter on Election Day https://t.co/R3ihQKTfvr
MLG__Will|GeorgeSulliho|0.296|0.0|0.82|0.18|@GeorgeSulliho gonna see how long I can join you with the election
sivanzustin|politico|0.6374|0.0|0.588|0.412|so trump is winning so far??? https://t.co/IoLyxD2sJx
infodude|ValaAfshar|0.0|0.0|1.0|0.0|RT @ValaAfshar: Past 10 election call times:1996: 9PM2000: December 12th2004: 11:19AM2008: 11PM20012: 11:17PM #ElectionNight https://
infodude||0.0|0.0|1.0|0.0|RT @ValaAfshar: Past 10 election call times:1996: 9PM2000: December 12th2004: 11:19AM2008: 11PM20012: 11:17PM #ElectionNight https://
niaimanix|JordinSparks|0.4559|0.094|0.684|0.222|"RT @JordinSparks: I'm praising the Lord right now! Because no matter what's happens in this election, HE STILL REIGNS! "
kvalandra2|bill_merkel|0.0|0.0|1.0|0.0|RT @bill_merkel: Media folk eat a helluva lot of pizza and cake on election days. At least according to all the photos I've seen today they
carolyncerbin|AmyBartner|0.0|0.0|1.0|0.0|RT @AmyBartner: We're broadcasting live on https://t.co/gLz3VscwjS with all your live election coverage! https://t.co/NJnVbC4SHZ
carolyncerbin|indystar|0.0|0.0|1.0|0.0|RT @AmyBartner: We're broadcasting live on https://t.co/gLz3VscwjS with all your live election coverage! https://t.co/NJnVbC4SHZ
PalatinateStyle|PalatinateUK|0.0|0.0|1.0|0.0|RT @PalatinateUK: Stay up to date with the latest from @PalatinatePoli1 as they cover the presidential race over night at: https://t.co/xBO
PalatinateStyle|t|0.0|0.0|1.0|0.0|RT @PalatinateUK: Stay up to date with the latest from @PalatinatePoli1 as they cover the presidential race over night at: https://t.co/xBO
ElectionGraphs|abulsme|0.0|0.0|1.0|0.0|VT/VA/GA/SC/IN/KY now closed. Only GA expected to be close. Others should be called relatively quickly. https://t.co/gmUwTGqJr4
JohnBahamonde1|MotherToEarthMV|0.0|0.0|1.0|0.0|RT @MotherToEarthMV: We are waiting for the election results to come it. https://t.co/WvQ0tGiIZ8
JohnBahamonde1|twitter|0.0|0.0|1.0|0.0|RT @MotherToEarthMV: We are waiting for the election results to come it. https://t.co/WvQ0tGiIZ8
K_rivera6|FriendlyAssh0le|0.8176|0.0|0.483|0.517|RT @FriendlyAssh0le: How I'm celebrating tonights election winner https://t.co/GKRWjQrEMQ
K_rivera6|twitter|0.8176|0.0|0.483|0.517|RT @FriendlyAssh0le: How I'm celebrating tonights election winner https://t.co/GKRWjQrEMQ
sleepingcolur|CNNPolitics|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
sleepingcolur|twitter|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
SocStudiesAPS|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
SocStudiesAPS|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
ford3102|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
EidojTrump|bunkerwsmith|0.5574|0.063|0.704|0.233|"RT @bunkerwsmith: To people feeling anxiety about the election: Focus on things you can control, like VOTING. Keep your chin up. Stay calm."
istx25|ughitsaaron|0.4767|0.0|0.78|0.22|RT @ughitsaaron: me &amp; my friends after this election is over https://t.co/D326G9pbVX
istx25|twitter|0.4767|0.0|0.78|0.22|RT @ughitsaaron: me &amp; my friends after this election is over https://t.co/D326G9pbVX
Ville_LNC|Cartel__shoota|0.0|0.0|1.0|0.0|"@Cartel__shoota @FearDept i dont think you can do ""right"" in this election"
Ligi20|CNN|0.25|0.0|0.895|0.105|"RT @CNN: Donald Trump peeked at Melania's ballot, and Twitter had some jokes. Big league. https://t.co/673JwvzlDn #ElectionDay https://t.co"
Ligi20|cnn|0.25|0.0|0.895|0.105|"RT @CNN: Donald Trump peeked at Melania's ballot, and Twitter had some jokes. Big league. https://t.co/673JwvzlDn #ElectionDay https://t.co"
MrMokelly|americanowradio|0.0|0.0|1.0|0.0|"RT @americanowradio: ELECTION 2016: What to watch for with @NikkiSchwab, @MrMokelly and @benfergusonshow HERE: https://t.co/BPxv2YIJTf http"
MrMokelly|americanowradio|0.0|0.0|1.0|0.0|"RT @americanowradio: ELECTION 2016: What to watch for with @NikkiSchwab, @MrMokelly and @benfergusonshow HERE: https://t.co/BPxv2YIJTf http"
1_Hit_Wonderful|Michaeljonair|0.5405|0.0|0.791|0.209|"RT @Michaeljonair: Not focused on #Election,can't stop thinking about hosting @BradPaisley on  #iHeartRadio Honda Stage LIVE This FRIDAY NI"
cesarcarvalho2|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
JohnWalsh001|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Movieguy2015|facebook|0.0|0.0|1.0|0.0|They left off the election process. Left off being qualified to run the country. https://t.co/wwLzq9s9Mu
ryan4moore99|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
SydneyyyAnn|POTUS|0.5093|0.0|0.68|0.32|"Favorite quote this election: ""Don't boo. Vote!"" - @POTUS"
ChrisDCBrau|oldglorybbq|0.4574|0.0|0.834|0.166|Find me upstairs on the patio at @oldglorybbq for The Corruption Election Party! #ElectionNight #voteogbbq https://t.co/0LxDwKOrlQ
ChrisDCBrau|twitter|0.4574|0.0|0.834|0.166|Find me upstairs on the patio at @oldglorybbq for The Corruption Election Party! #ElectionNight #voteogbbq https://t.co/0LxDwKOrlQ
Karoli|cmwarnerstl|0.0|0.0|1.0|0.0|@cmwarnerstl we have a live blog going here! https://t.co/WUWaqEdKxG
Karoli|crooksandliars|0.0|0.0|1.0|0.0|@cmwarnerstl we have a live blog going here! https://t.co/WUWaqEdKxG
JB93621|GoAngelo|0.0|0.0|1.0|0.0|"RT @GoAngelo: Election Night 2012Actual ResultsObama: 65,915,795Romney: 60,933,504 https://t.co/dtD8WwpAd6"
JB93621|twitter|0.0|0.0|1.0|0.0|"RT @GoAngelo: Election Night 2012Actual ResultsObama: 65,915,795Romney: 60,933,504 https://t.co/dtD8WwpAd6"
marcooviedo|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
marcooviedo|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
AndrewGilbert1|InTheSoupAgain|0.7772|0.0|0.658|0.342|"RT @InTheSoupAgain: Listening to @BBCRadio4 election new special. Rather good, not as depressing as I thought it would be."
WallyWaffles27|JeremyMcLellan|0.5423|0.079|0.717|0.204|RT @JeremyMcLellan: There is no greater testament to the strength of the Muslim community than that they made it through this election with
bjohnsmeyer|jodyavirgan|-0.431|0.185|0.815|0.0|@jodyavirgan your wit is getting me through this election. Don't listen to the people that don't like dad jokes.
schorpp1955|msn|0.0|0.0|1.0|0.0|Election 2016 https://t.co/lap23s1KrR
unfilunfet|JohnKingCNN|0.0|0.0|1.0|0.0|@JohnKingCNN in mid election season form on the board tonight! Make that board sing John. #hemaybeawizard  #Election2016 #ElectionNight
Tjudge34|Robertzul2|0.5719|0.0|0.812|0.188|@Robertzul2 If trumo wins the election this country is screwed.....  He's a dictator......  Impeached in less than a year
LexiLips|Things4WhitePpl|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
LexiLips|twitter|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
scr385w|NRO|0.0|0.0|1.0|0.0|"RT @NRO: Early Exit Polls: Trump Opens YUGE Gap between College-Educated, Non-College-Educated Whiteshttps://t.co/ADpCNhYfiC #ElectionNight"
kayleenkrafft|EbingerTrey|-0.2782|0.141|0.759|0.1|RT @EbingerTrey: So whose ready for war with Russia? Cause depending on the way this election is leaning we will be having a draft
WmScottBlair|FeliciaBGomez|-0.298|0.149|0.744|0.106|"RT @FeliciaBGomez: Translation: ""We just realized that Hillary's LOSING in NC! Quick! Change the rules! Who cares if it's on the actual ele"
gravity_jo|twitter|0.101|0.0|0.878|0.122|Election Day today. Vote for the stuff that fucking matters https://t.co/6E28hDjkeJ
CammStride|foxnews|0.0|0.0|1.0|0.0|"Here's my prediction. What do ya think, fellow centipedes?? #Election2016 #ElectionNight #MAGA #MAGA3x https://t.co/0LSZB7OBaP"
muppetaphrodite|WaltDisneyWorld's|0.0|0.0|1.0|0.0|Election night escapism at @WaltDisneyWorld's Sanaa. https://t.co/10ZlQTUz02
muppetaphrodite|twitter|0.0|0.0|1.0|0.0|Election night escapism at @WaltDisneyWorld's Sanaa. https://t.co/10ZlQTUz02
waughbr|seanhannity|0.0|0.0|1.0|0.0|@seanhannity @realDonaldTrump frank lungs just called the election for Hillary?
nathanbship|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
nathanbship|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
lavventuras|Maddynx|0.0|0.0|1.0|0.0|RT @Maddynx: Twitter on Election Dayhttps://t.co/04p0nkjyiw
Gustavwasa1|twitter|0.5719|0.0|0.709|0.291|Happy Election Day to the voters &amp; volunteers everywhere. https://t.co/qkEENOed4I
hughmooney1|artfinder|0.0|0.0|1.0|0.0|ARTFINDER: US Election night by Hugh Mooney - Acrylic paint and  polystyrene skull on found c... - https://t.co/YQVOf1B6EK via @artfinder
hughmooney1|artfinder|0.0|0.0|1.0|0.0|ARTFINDER: US Election night by Hugh Mooney - Acrylic paint and  polystyrene skull on found c... - https://t.co/YQVOf1B6EK via @artfinder
caroletalk|WDFx2EU8|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
caroletalk|conservativeeagles|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
vgc120|JonErlichman|0.0|0.0|1.0|0.0|RT @JonErlichman: Things that didn't exist election night in 2008:UberiPadInstagramSnapchatWhatsAppPinterestPeriscopeOculusSlack
kshwiff|WSJPolitics|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
kshwiff|wsj|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
gocoo|LanceBass|0.0|0.0|1.0|0.0|RT @LanceBass: Lily's first election dingofosterlily #ElectionDay #ImWithHer https://t.co/myazwZQb7P
gocoo|instagram|0.0|0.0|1.0|0.0|RT @LanceBass: Lily's first election dingofosterlily #ElectionDay #ImWithHer https://t.co/myazwZQb7P
Kinniska|SamuraiKnitter|-0.2732|0.213|0.667|0.12|"@SamuraiKnitter and yes, I'm hiding in pedantry as a distraction from the election. Less heartburn than alcohol this way."
journobeth|nymag|0.0|0.0|1.0|0.0|"If this race *is* settled early, we can all turn our focus to the less nerve-wracking, more entertai ..  https://t.co/FSTure4CR2"
Dinahmente|LaurenJauregui|0.4795|0.0|0.881|0.119|RT @LaurenJauregui: I'm so excited that I was able to exercise my vote as a Cuban American Woman for the first time in this particular elec
karymeolivera_9|callliiee__|-0.5267|0.348|0.489|0.163|RT @callliiee__: This election got everyone hating each other. It's honestly sad
JJ7701|SueCFlorida|-0.1531|0.068|0.932|0.0|"RT @SueCFlorida: For the first time in 20 years, I will not be watching @FoxNews Election Coverage. I can't stand Megyn Kelly. Will miss @B"
997wtn|WildWingCafeTN|0.4574|0.0|0.864|0.136|Our stage is set! We're about 30 mins away from broadcasting live at @WildWingCafeTN for this year's Election Party https://t.co/G2ceN9Llil
997wtn|twitter|0.4574|0.0|0.864|0.136|Our stage is set! We're about 30 mins away from broadcasting live at @WildWingCafeTN for this year's Election Party https://t.co/G2ceN9Llil
Gunning_96|NHL|0.3818|0.0|0.843|0.157|RT @NHL: On this Election Day there is only one clear choice. #ImWithPhil #MakeAmericaSkateAgain https://t.co/DXGnvMX1Of
Gunning_96|twitter|0.3818|0.0|0.843|0.157|RT @NHL: On this Election Day there is only one clear choice. #ImWithPhil #MakeAmericaSkateAgain https://t.co/DXGnvMX1Of
Noodlepig|FOXnews2016|0.6801|0.0|0.682|0.318|@FOXnews2016  In U.K. Watching the election. Most importantly show us the 'Sweet Shorts'. #FoxNews2016
BroadNOLA|us9|-0.1984|0.218|0.635|0.147|Happy Election Day! Forget your troubles with a quick read of our newsletter. We open ARRIVAL &amp; CHRISTINE on Friday!https://t.co/tFMs0hd2am
TheTekFanatic|Trump2016Pence|-0.8979|0.459|0.541|0.0|"RT @Trump2016Pence: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
TheTekFanatic||-0.8979|0.459|0.541|0.0|"RT @Trump2016Pence: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
Minimaria|AJEnglish|0.0|0.0|1.0|0.0|RT @AJEnglish: Here's when to expect election results.Follow the live results here: https://t.co/arXvIMQVja #ElectiondDay #Election2016 ht
Minimaria|interactive|0.0|0.0|1.0|0.0|RT @AJEnglish: Here's when to expect election results.Follow the live results here: https://t.co/arXvIMQVja #ElectiondDay #Election2016 ht
AdedigbaAdeniy1|washingtonpost|0.3612|0.0|0.839|0.161|"RT @washingtonpost: A Trump presidency would be like Stevie Wonder driving, Stevie Wonder says https://t.co/tLNfxuxYPc"
AdedigbaAdeniy1|washingtonpost|0.3612|0.0|0.839|0.161|"RT @washingtonpost: A Trump presidency would be like Stevie Wonder driving, Stevie Wonder says https://t.co/tLNfxuxYPc"
SuadAbdalla44|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
SuadAbdalla44|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
RyanWoodDFW|wusa9!|0.0|0.0|1.0|0.0|Election night at @wusa9!  @joanievas and I are heading up central coverage for @TEGNA!  
alice__baek|JackHoward|0.0|0.0|1.0|0.0|RT @JackHoward: I can't vote in this election but if I could I would vote for the first woman president after the first black president. Be
poe_slilraven|instagram|0.8346|0.0|0.67|0.33|Thank you Aunt Carla for taking me to vote in my first election!! You're the best!! #noexcuses https://t.co/f8djt1TTpE
captainamarigan|dacthe2|-0.7351|0.437|0.563|0.0|RT @dacthe2: Sick and tired of hearing about this election
Brrend99|zachhaller|-0.4215|0.118|0.882|0.0|RT @zachhaller: Shed a tear when I found out my sister #voted @DrJillStein in her 5th grade mock electionJill earned my vote tooThis 1's
BrianLockwood|MNN59|-0.079|0.204|0.612|0.184|"liking @MNN59 live coverage of the election, feels less stressful https://t.co/7iY609QiXt"
BrianLockwood|livestream|-0.079|0.204|0.612|0.184|"liking @MNN59 live coverage of the election, feels less stressful https://t.co/7iY609QiXt"
serena_223|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
serena_223|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
Alan_Sky|twitter|0.0|0.0|1.0|0.0|Holy cow! This ad during US election night...  https://t.co/ArgPyCHOwz
nikipressey77_p|IMIXWHATILIKE|0.296|0.0|0.901|0.099|RT @IMIXWHATILIKE: I voted for @DrJillStein - Join me and @ajamubaraka and others tonight at 7p EST for our election night coverage  https:
DJseancurtisJNR|andrewismaxwell|0.0|0.0|1.0|0.0|"RT @andrewismaxwell: So here we go,polls closing..The very first U.S. election between a candidate and a contestant.#ElectionNight"
hcollis|politico|-0.1531|0.118|0.882|0.0|Follow #election day liveblog with POLITICO including the 16 battlegrounds to watch: https://t.co/6mI5M1IFOh
JohnRClem|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
ChrissyFisch_PF|RickMitchellWX|0.0|0.0|1.0|0.0|RT @RickMitchellWX: Fueling up for a busy night of election coverage. #nbcdfw https://t.co/fRok4sVbsN
ChrissyFisch_PF|twitter|0.0|0.0|1.0|0.0|RT @RickMitchellWX: Fueling up for a busy night of election coverage. #nbcdfw https://t.co/fRok4sVbsN
webandgraphix|digitaltrends|0.3818|0.0|0.809|0.191|Electionland Google Trends map helps voters visualize polling station issues https://t.co/x9TqzPcDDa https://t.co/6Q1P8f8orL
rollx3|nprpolitics|0.0|0.0|1.0|0.0|"RT @nprpolitics: For full coverage and analysis, follow our live blog. https://t.co/0WfRXoXnye #ElectionDay #Election2016 https://t.co/Rcqe"
rollx3|npr|0.0|0.0|1.0|0.0|"RT @nprpolitics: For full coverage and analysis, follow our live blog. https://t.co/0WfRXoXnye #ElectionDay #Election2016 https://t.co/Rcqe"
RiannaTweeet|WorkingBarbie|-0.6597|0.229|0.706|0.065|"RT @WorkingBarbie: Waiting for election results is like waiting for a grade on a group project. I know I did my shit right, but I'm scared"
EastBayTimes|eastbaytimes|0.0|0.0|1.0|0.0|Election Night live blog: Results and updates https://t.co/r4uWNieZ9E https://t.co/1xVwme9iJN
steelrsfan57|katehansen21|0.6115|0.0|0.79|0.21|RT @katehansen21: it's the most wonderful time of the year (#Election Day) #ImWithHer #Election2016 #OHHillYes https://t.co/JY4Hm6jKhJ
steelrsfan57|twitter|0.6115|0.0|0.79|0.21|RT @katehansen21: it's the most wonderful time of the year (#Election Day) #ImWithHer #Election2016 #OHHillYes https://t.co/JY4Hm6jKhJ
ideavator|FreddieCampion|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
ideavator|twitter|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
Navyboy08021|MaryLoveUS4|0.0|0.0|1.0|0.0|RT @MaryLoveUS4: BREAKING: All Election Systems Are Down in Swing State of Colorado https://t.co/j3TKvwf6lS https://t.co/WtCJ1yHL1r
Navyboy08021|conservativetribune|0.0|0.0|1.0|0.0|RT @MaryLoveUS4: BREAKING: All Election Systems Are Down in Swing State of Colorado https://t.co/j3TKvwf6lS https://t.co/WtCJ1yHL1r
SueCFlorida|FredZeppelin12|0.25|0.0|0.895|0.105|RT @FredZeppelin12: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERS. Advantage #Trump. Evening voters are evening voters because t
VogueRunway|vogue|0.5777|0.0|0.681|0.319|Doing your civic duty never looked so good. https://t.co/3mUf48wbzc
Khaleesi_Hodan|TheDailyShow|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
Khaleesi_Hodan|cc|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
hunterlurie|SeanMBurns|0.2023|0.0|0.909|0.091|@SeanMBurns @mattzollerseitz it's important that the price tag for his screenplay about this year's election be at least $10M
syed_allauddin|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
syed_allauddin|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
AnisaGohar|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
AnisaGohar|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
sagegoharirfan1|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
sagegoharirfan1|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
IrfanGohar02|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
IrfanGohar02|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
mfiusa01|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
mfiusa01|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
JayDizL04|lolrenaynay|0.4939|0.086|0.703|0.211|"RT @lolrenaynay: Election results come in soon, come here and let me save youFYI I'm drinkingYou can join me, no judgementhttps://t.co/S"
IrfanGohar4|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
IrfanGohar4|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
dangerdan8|Ls_Up_850|0.0|0.0|1.0|0.0|RT @Ls_Up_850: NSD &gt; President election Location on if you wanna debate physically
Anisairfan2|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
Anisairfan2|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
crewelladevil|ChristnHipster|0.0|0.0|1.0|0.0|RT @ChristnHipster: what to do instead of watching election coverageread dostoevskylisten to sufjansmoke a pipefinger paintsip a stou
IrfanGohar|mehdifoundation|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
IrfanGohar|medium|0.0|0.0|1.0|0.0|RT @mehdifoundation: #Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNig
KingKinthehouse|TeenVogue|-0.3595|0.333|0.667|0.0|"RT @TeenVogue: No peeking, Donald! https://t.co/Q2GflxtECB"
KingKinthehouse|teenvogue|-0.3595|0.333|0.667|0.0|"RT @TeenVogue: No peeking, Donald! https://t.co/Q2GflxtECB"
chrissyrules66|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
miyuwi|CNN|0.0|0.0|1.0|0.0|RT @CNN: This is how close Clinton and Trump will be to each other in Manhattan tonight https://t.co/YPAfWQsye5 #ElectionDay https://t.co/4
miyuwi|cnn|0.0|0.0|1.0|0.0|RT @CNN: This is how close Clinton and Trump will be to each other in Manhattan tonight https://t.co/YPAfWQsye5 #ElectionDay https://t.co/4
KB_v3|twitter|0.0|0.0|1.0|0.0|"Election Day is the day that the nation disobeys s national rule, talking about politics https://t.co/Y6x0HzhyQa"
joelbthomas|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
joelbthomas|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
StephanieMitz|FemMajority|0.0|0.0|1.0|0.0|"RT @FemMajority: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https"
TuNaLdO|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
TuNaLdO|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
piquergaming|twitter|0.0|0.0|1.0|0.0|Updating my Election Day soundtrack: https://t.co/MjDnNKSpYA
bryanclark|twitter|0.0|0.0|1.0|0.0|BuzzFeed's live election coverage is 'Ow My Balls' IRL #ElectionNight https://t.co/l8NcxeHyN2
GalloCostantino|AaronBlake|0.0|0.0|1.0|0.0|RT @AaronBlake: 8 states that will tell you everything you need to know on tonight https://t.co/Q3yZLpiufZ https://t.co/t5mguPjnGv
GalloCostantino|washingtonpost|0.0|0.0|1.0|0.0|RT @AaronBlake: 8 states that will tell you everything you need to know on tonight https://t.co/Q3yZLpiufZ https://t.co/t5mguPjnGv
BrandConverts|SebGorka|0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
BrandConverts||0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
DouglasRojas|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
DouglasRojas|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
dmarieolsen|bpmoritz|0.0|0.0|1.0|0.0|RT @bpmoritz: Pizza is filtering into newsrooms around the country. Eyes are rolling in adjacent sports departments. https://t.co/60ORNPGmfy
dmarieolsen|sportsmediaguy|0.0|0.0|1.0|0.0|RT @bpmoritz: Pizza is filtering into newsrooms around the country. Eyes are rolling in adjacent sports departments. https://t.co/60ORNPGmfy
BaileeBolt|MattMoretta|0.8934|0.0|0.545|0.455|"RT @MattMoretta: Plot twist: Matthew McConaughey wins election, everyone receives a brand new Lincoln, happiness is restored alright alrigh"
ShainEThomas|CNN|0.0|0.0|1.0|0.0|"""Stand by for projection"" https://t.co/gV2CluIl9U via @CNN"
ShainEThomas|linkis|0.0|0.0|1.0|0.0|"""Stand by for projection"" https://t.co/gV2CluIl9U via @CNN"
Dowling_Sam|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
complex_roolz|theverge|0.0|0.0|1.0|0.0|Status Update: 10 provocative political novels to read after the election https://t.co/Wv9PmoxmfU
edward_thefirst|DavMicRot|0.7579|0.0|0.755|0.245|"RT @DavMicRot: Clinton up to 91% #President on strength of strong turnout in Florida which is up to 87% https://t.co/kZWGoxX4EF slow, stead"
edward_thefirst|predictwise|0.7579|0.0|0.755|0.245|"RT @DavMicRot: Clinton up to 91% #President on strength of strong turnout in Florida which is up to 87% https://t.co/kZWGoxX4EF slow, stead"
drmojo1975|ArcticFox2016|-0.5904|0.215|0.785|0.0|RT @ArcticFox2016: PROOF That Censorship Against Conservatives is WORSE as Election Day Approaches [Video] https://t.co/PQJmVRONI0
drmojo1975|conservativevideos|-0.5904|0.215|0.785|0.0|RT @ArcticFox2016: PROOF That Censorship Against Conservatives is WORSE as Election Day Approaches [Video] https://t.co/PQJmVRONI0
brianaaaxMH|SheHatesJacoby|0.5719|0.0|0.748|0.252|RT @SheHatesJacoby: Back in 2012 when Obama won the 2012 election https://t.co/QgQ76yrR2l
brianaaaxMH|twitter|0.5719|0.0|0.748|0.252|RT @SheHatesJacoby: Back in 2012 when Obama won the 2012 election https://t.co/QgQ76yrR2l
Jaredddd123|Capitals|0.0|0.0|1.0|0.0|RT @Capitals: The #Gr8 has spoken. #VoteWilson Follow #CapsElectionNight results: https://t.co/NaZbAPTUBj https://t.co/Q6VoebJap3
Jaredddd123|nhl|0.0|0.0|1.0|0.0|RT @Capitals: The #Gr8 has spoken. #VoteWilson Follow #CapsElectionNight results: https://t.co/NaZbAPTUBj https://t.co/Q6VoebJap3
politicallyrich|RT_America|0.0|0.0|1.0|0.0|RT @RT_America: BREAKING: WikiLeaks releases election day batch from Clinton campaign chair #podestaemails35 https://t.co/gvkGurkYr9 https:
politicallyrich|rt|0.0|0.0|1.0|0.0|RT @RT_America: BREAKING: WikiLeaks releases election day batch from Clinton campaign chair #podestaemails35 https://t.co/gvkGurkYr9 https:
hotteronline|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
barbya1|slone|0.0|0.0|1.0|0.0|"RT @slone: ELECTION WILL BE DECIDED BY EVENING VOTERS**PROJECTED 140 MILLION TOTAL**SHOWDOWN: FL, MI, NC, PAhttps://t.co/hb7QtnFCiq"
TWEETY021163|globeandmail|-0.4019|0.153|0.847|0.0|RT @globeandmail: America votes: Polls in some battleground states set to close soon https://t.co/9CWjksdux4 #ElectionNight #Election2016
TWEETY021163|theglobeandmail|-0.4019|0.153|0.847|0.0|RT @globeandmail: America votes: Polls in some battleground states set to close soon https://t.co/9CWjksdux4 #ElectionNight #Election2016
ChadAinsworth|instagram|0.0|0.0|1.0|0.0|Watching the election results tonight as a family with a little Caps https://t.co/k5lkvDLlVA
News__La|CBSNews|0.2716|0.0|0.909|0.091|RT @CBSNews: First exit poll of Election 2016 shows that the most important issue to North Carolina is the economy #Election2016 https://t.
News__La||0.2716|0.0|0.909|0.091|RT @CBSNews: First exit poll of Election 2016 shows that the most important issue to North Carolina is the economy #Election2016 https://t.
marjoriemliu|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
marjoriemliu|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
Vi_Cos|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
Vi_Cos|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
JoeLeydon|Glenn__Kenny|-0.4005|0.109|0.891|0.0|@Glenn__Kenny Wife &amp; I went to see Marty Robbins perform on Election Day 80 - after networks called it for Reagan. We got very drunk.
bolajoselopez|JordanHyland21|0.3182|0.103|0.7|0.198|RT @JordanHyland21: If Donald Trump wins the election I will Paypal $100 to one person who retweets this. No backing out.
AguiRuben|SoaRPraizist|0.5719|0.0|0.802|0.198|"RT @SoaRPraizist: If Trump wins the election, I will make artwork for everyone that RTs this tweet"
HaroMariana|THR|0.6369|0.0|0.625|0.375|RT @THR: Hollywood's best #Election2016 tweets https://t.co/FJx6s6ouYO https://t.co/PmPwzeyzE4
HaroMariana|hollywoodreporter|0.6369|0.0|0.625|0.375|RT @THR: Hollywood's best #Election2016 tweets https://t.co/FJx6s6ouYO https://t.co/PmPwzeyzE4
ElxseM|triIIfenty|0.296|0.0|0.761|0.239|RT @triIIfenty: This whole election is a joke https://t.co/OZrOXX7iFJ
ElxseM|twitter|0.296|0.0|0.761|0.239|RT @triIIfenty: This whole election is a joke https://t.co/OZrOXX7iFJ
tomthelitgeek|uniofeastanglia|0.2732|0.115|0.718|0.167|In media centre preparing for election shift 1.30am https://t.co/GqUhH0c3tf as @uniofeastanglia gone crazy tonight... gonna be fascinating
tomthelitgeek|livewire1350|0.2732|0.115|0.718|0.167|In media centre preparing for election shift 1.30am https://t.co/GqUhH0c3tf as @uniofeastanglia gone crazy tonight... gonna be fascinating
GreenBiotechie|chrislhayes|-0.5256|0.159|0.841|0.0|RT @chrislhayes: Trump is already laying the groundwork to contest the legitimacy of the election and it's incredibly dangerous.
Nikki_Bitchhh|ShineVista|0.3616|0.148|0.608|0.243|"RT @ShineVista: Prediction: Hillary Clinton wins election, Donald Trump doesn't concede. America riots, &amp; people die. Market crashes. Haram"
Saritrovick|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
Saritrovick|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
tracieabrennan|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
HandballGardien|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
HandballGardien|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
eliglazier|Devon2012|-0.1779|0.086|0.914|0.0|"@Devon2012 seriously. this fucking guy doesnt TELL ANYONE who hes voting for until 6:30pm on Election Day, the schmuck."
joeybaker09|RealJeremyNolt|-0.6124|0.238|0.762|0.0|"RT @RealJeremyNolt: CNN: Rigged a debate, rigged interviews, colluded with the DNC, then told everyone the election wasn't rigged.#MAGA#"
scarpetta70|hardball|0.6369|0.0|0.781|0.219|RT @hardball: I personally think its the best part of politics  the concession speech. -- @HardballChris https://t.co/Fsziwkk70U
scarpetta70|variety|0.6369|0.0|0.781|0.219|RT @hardball: I personally think its the best part of politics  the concession speech. -- @HardballChris https://t.co/Fsziwkk70U
Mangoluu|crooksandliars|0.6996|0.0|0.674|0.326|RT @crooksandliars: Join @Karoli and the whole @crooksandliars crew for Election night fun! https://t.co/wee0H8Tgb7
Mangoluu|crooksandliars|0.6996|0.0|0.674|0.326|RT @crooksandliars: Join @Karoli and the whole @crooksandliars crew for Election night fun! https://t.co/wee0H8Tgb7
ranakhalifeh|chrisbharrison|0.0|0.0|1.0|0.0|RT @chrisbharrison: Tonight..in the most dramatic election ever..2 candidates..only one will make it to the White House (read in Harrison v
AdamInBako|WalshFreedom|-0.4019|0.351|0.649|0.0|RT @WalshFreedom: Who gives a damn? https://t.co/rJWutS0KlH
AdamInBako|thehill|-0.4019|0.351|0.649|0.0|RT @WalshFreedom: Who gives a damn? https://t.co/rJWutS0KlH
Rempancy|abittoolethal|0.0|0.0|1.0|0.0|RT @abittoolethal: LIVEPracticing for post-2016 Presidential election || #TheDivision Survivalhttps://t.co/D94UmH7JOw
Gamer2012Pro|ReutersPolitics|0.0|0.0|1.0|0.0|RT @ReutersPolitics: Factbox: State-by-state poll closing times for U.S. election https://t.co/KW4DXXwRK0 https://t.co/A0GOWkdonw
Gamer2012Pro|reuters|0.0|0.0|1.0|0.0|RT @ReutersPolitics: Factbox: State-by-state poll closing times for U.S. election https://t.co/KW4DXXwRK0 https://t.co/A0GOWkdonw
_onlyonequeen|HaleeSharp13|0.4877|0.0|0.869|0.131|RT @HaleeSharp13: The only thing this election has shown me is that Jesus is coming back very soon. Y'all better start prayin' 
patriciayingst|WSJ|-0.4767|0.162|0.838|0.0|RT @WSJ: An online attack disrupted call operations for Clintons presidential campaign ahead of Tuesdays election https://t.co/aOAAprwBob
patriciayingst|wsj|-0.4767|0.162|0.838|0.0|RT @WSJ: An online attack disrupted call operations for Clintons presidential campaign ahead of Tuesdays election https://t.co/aOAAprwBob
GregIenco|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
GregIenco|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
DoloresWells20|WSJPolitics|0.0|0.0|1.0|0.0|"RT @WSJPolitics: At 7 p.m., polls close in six states, including some that could signal where this race is headed. Live analysis: https://t"
DoloresWells20||0.0|0.0|1.0|0.0|"RT @WSJPolitics: At 7 p.m., polls close in six states, including some that could signal where this race is headed. Live analysis: https://t"
TeresaE17|hrtablaze|0.9207|0.0|0.645|0.355|RT @hrtablaze: My Bernie Sanders loving nephew who has been messing with me all election just told me he voted TRUMP !!! WOOT WOOT ! #elect
OJkimson|jessesingal|0.6369|0.0|0.741|0.259|"RT @jessesingal: Single best video clip of Election Day so far, hands downhttps://t.co/uiPEsSdkIp"
andyparmo|FrizFrizzle|-0.7096|0.237|0.763|0.0|RT @FrizFrizzle: MOVIE IDEA: Lightning strikes the BBC on Election Night and Jeremy Vine is trapped in his CGI Results World.
klintevans|Wu_Tang_Finance|0.0|0.0|1.0|0.0|RT @Wu_Tang_Finance: The 2016 election we deserve https://t.co/7uY6L705xS
klintevans|twitter|0.0|0.0|1.0|0.0|RT @Wu_Tang_Finance: The 2016 election we deserve https://t.co/7uY6L705xS
jamesdouglasm11|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
RobertsBumbaugh|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
RobertsBumbaugh|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
BComp272|WSJPolitics|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
BComp272|wsj|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
UsmanUmar199|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
UsmanUmar199|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
WorldOfStu|lostfreak4|0.7612|0.0|0.681|0.319|"@lostfreak4 I mean yes, but its election day so I force my hand.  Put it in the D column."
Littleone619|bfraser747|0.0|0.0|1.0|0.0|RT @bfraser747:  #NeverHillaryThis election isn't about Rep vs. Dem. It's about #Corruption vs #MAGA#Election2016 #VoteTrump#Electi
yoAfrodite|twitter|0.7645|0.0|0.548|0.452|I wish I had more positive feelings about this election but... https://t.co/Ilg4cl0ej6
_solleb|FreddieCampion|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
_solleb|twitter|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
BeyNa_PalyNa|Nigel_Farage|0.4767|0.051|0.809|0.14|RT @Nigel_Farage: Enjoyed speaking to @Varneyco earlier. @realDonaldTrump represents change in this election just as Leave did in the EU re
JJP1952|twitter|-0.0772|0.124|0.769|0.107|MSNBC is on top of this election. I wonder why their ratings are always low? https://t.co/DXTfZvf58h
KayHillYes|Emory4Hillary|0.0|0.0|1.0|0.0|"RT @Emory4Hillary: BREAKING NEWS: Election Update, some precincts in Georgia will remain open until 7:30 pm due to high voter turnout. Keep"
Morgan_Rawlss|kurtsteiss|0.0|0.0|1.0|0.0|"RT @kurtsteiss: There are now 6,884 flags on the #okstate library lawn, and they aren't for the election. Each flag represents a soldier ki"
KBDanquah|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
KBDanquah|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
LMSNCUS|DrMartyFox|-0.0173|0.131|0.741|0.128|RT @DrMartyFox: This Election Is NOT A Choice Between The Lesser Of Two Evils This Is A Choice Between GOOD &amp; PURE EVIL#Voted #Trump On
Lope_Doggg|jerm_rice|-0.34|0.146|0.854|0.0|RT @jerm_rice: There's gonna be a fire movie/series about this election a few years down the road
osnapitsjoyce|KathleenLights1|0.4199|0.141|0.573|0.286|RT @KathleenLights1: Hope everyone voted today! This election has traumatized me.... I pray for America.
imscottmorris|twitter|0.4939|0.0|0.652|0.348|This election's pretty much done... #vote2016 https://t.co/cCxlLu3ehI
Adeline_Garrett|YURlPlRATE|0.6633|0.0|0.783|0.217|RT @YURlPlRATE: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
FiveThirtyEight|fivethirtyeight|0.0|0.0|1.0|0.0|The people elected today will affect when (if??) we get to Mars. #ElectionNight https://t.co/CbMh5dTJ0E https://t.co/PaD0DzxyM0
stirlospace|_alastair|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
stirlospace|t|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
hannahxalicea|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
G_Stratt|barstoolsports|0.5719|0.0|0.856|0.144|"RT @barstoolsports: Before you move to Canada after this election, learn some more about our neighbors to the north. They're happy to have"
jwinks_17|SavageBoySoy|0.0|0.0|1.0|0.0|RT @SavageBoySoy: After tonight's election https://t.co/gkakonQZKz
jwinks_17|twitter|0.0|0.0|1.0|0.0|RT @SavageBoySoy: After tonight's election https://t.co/gkakonQZKz
panicstlawyer|ESPNStatsInfo|0.34|0.0|0.906|0.094|RT @ESPNStatsInfo: Connor McDavid &amp; Sidney Crosby meet for 1st timeMario Lemieux &amp; Wayne Gretzky played vs each other for 1st time on Ele
Namndhela|Seantaneous|0.0|0.0|1.0|0.0|RT @Seantaneous: it is now election day. https://t.co/olmaUaOnC9
Namndhela|twitter|0.0|0.0|1.0|0.0|RT @Seantaneous: it is now election day. https://t.co/olmaUaOnC9
Caarmsssss|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
CCrusherP|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
camilabellenn|Arianaajpg|-0.6124|0.211|0.789|0.0|RT @Arianaajpg: this election has brought out all the racist people that still exist in America...sad
Thetenorplayer|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
Thetenorplayer|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
pinkkstarbucks|CNN|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
pinkkstarbucks|twitter|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
alisonrose711|voxdotcom|0.0|0.0|1.0|0.0|RT @voxdotcom: #MyMuslimVote lets Muslims speak for themselves  finally https://t.co/3ySZq9p54T
alisonrose711|vox|0.0|0.0|1.0|0.0|RT @voxdotcom: #MyMuslimVote lets Muslims speak for themselves  finally https://t.co/3ySZq9p54T
jadanicolexo_|ynrichards|0.0|0.0|1.0|0.0|RT @ynrichards: Election Day is NOT Inauguration DayElection Day is NOT Inauguration DayElection Day is NOT Inauguration DayElection Day
Politicianist|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
Politicianist|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
KickinItWithKae|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
KickinItWithKae|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
amandaberkshire|annehelen|-0.1645|0.111|0.8|0.089|RT @annehelen: the piece I've been writing in my head all year &amp; my last of the election cycle: Don't Cry for Ivanka Fear Herhttps://t.
murphyj21|surfermom77|0.0|0.0|1.0|0.0|"RT @surfermom77: Twitter &amp; FB R begin inundated wt reports of Elec.fraud, voting irregularities &amp; discrimination against Trump Votershttps"
fruace|oneofonealbum|0.5719|0.0|0.821|0.179|RT @oneofonealbum: If Trump   Wins The Election I Am Moving   Out Of The Country  Goodbye   America   Hello   SHINee Wo
WagnerJwagner23|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
pg_countryboy|LifeAsRednecks|0.0|0.0|1.0|0.0|RT @LifeAsRednecks: Election Prediction: Democrats take an early lead until Republicans finally get off work to go and vote
DonaldTrumpNewz|endingthefed|-0.5319|0.278|0.605|0.118|"URGENT  George Soros Secret Plot to STEAL Election Has Been EXPOSED, Spread This Around https://t.co/uByA63hei8 https://t.co/32enxEBGEh"
HerbApproach|theweedblog|0.0|0.0|1.0|0.0|Why Hillary Clinton Could be More Than the First https://t.co/22pBl7AV3J #Ending_Marijuana_Prohibition #election_2016 #hillary_clinton
_Scyx|PeIicans|0.0|0.0|1.0|0.0|RT @PeIicans: Election prediction: Democrats to take an early lead which will change once Republicans get off work and are able to vote.
mbuckbee|joeyalison|-0.8779|0.336|0.664|0.0|"RT @joeyalison: Me just now: Oh, fuck, what the fuck is this election map, oh jesus...wait, this is a goddamn cell phone ad. https://t.co/h"
mbuckbee|t|-0.8779|0.336|0.664|0.0|"RT @joeyalison: Me just now: Oh, fuck, what the fuck is this election map, oh jesus...wait, this is a goddamn cell phone ad. https://t.co/h"
DoctorBuxter|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
FACT_gr|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
FACT_gr|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
CoreyRYung|fivethirtyeight|0.2023|0.0|0.899|0.101|How important is Florida? (Polls in the eastern part of the stateclose in a few minutes.) If https://t.co/c42reO6IbC
MCRWillCarryOn_|BoofBaldy|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
MCRWillCarryOn_|twitter|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
dale_bernadette|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
dale_bernadette||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
ColleenChaaland|ransom54|-0.5927|0.188|0.812|0.0|RT @ransom54: Already did. Will boycott them after the election too. I don't have any desire to return to those networks at all! https://t.
ColleenChaaland||-0.5927|0.188|0.812|0.0|RT @ransom54: Already did. Will boycott them after the election too. I don't have any desire to return to those networks at all! https://t.
jansims471|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
bresenpai|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
bresenpai|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
iYousif|AnsonWhaley|0.0|0.0|1.0|0.0|RT @AnsonWhaley: This is absolutely the only way the first vote could have been registered in this election. https://t.co/qhoJ4AJe0q
iYousif|vine|0.0|0.0|1.0|0.0|RT @AnsonWhaley: This is absolutely the only way the first vote could have been registered in this election. https://t.co/qhoJ4AJe0q
election_votes|scaryycsgo|0.0|0.0|1.0|0.0|RT @scaryycsgo: Who are you voting for this election? #ElectionNight #electionday #ElectionFinalThoughts
issa_abutaa|ajplus|0.636|0.0|0.819|0.181|"RT @ajplus: We're loving the 'I VOTED' selfies and #ElectionDay stories you're sending our FB Messenger election bot, Mila! https://t.co/QQ"
issa_abutaa|t|0.636|0.0|0.819|0.181|"RT @ajplus: We're loving the 'I VOTED' selfies and #ElectionDay stories you're sending our FB Messenger election bot, Mila! https://t.co/QQ"
mariapaularomo|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
mariapaularomo|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
lisadunny40|itvnews|0.0|0.0|1.0|0.0|"RT @itvnews: Follow ITV News' election night coverage live on Facebook, or tune in to ITV from 10.40pmhttps://t.co/rplwx2DhfI #Election201"
Daniso|WSJ|0.5719|0.0|0.837|0.163|"RT @WSJ: Obama isnt on the ballot, but early exit-poll results show he's popular among the U.S. electorate https://t.co/XFnrzvuItF  #Elec"
Daniso|wsj|0.5719|0.0|0.837|0.163|"RT @WSJ: Obama isnt on the ballot, but early exit-poll results show he's popular among the U.S. electorate https://t.co/XFnrzvuItF  #Elec"
LilyDirection7|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
LilyDirection7|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
AdvHoustonChiro|portacle|0.7065|0.0|0.405|0.595|This Election - SHARE SHARE SHARE|Portacle https://t.co/LNKwPkb0gZ
chelseabowen|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
chelseabowen|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
AaronBastani|novaramedia|0.0|0.0|1.0|0.0|My people tell me I'll be here all night https://t.co/LhaB86IEcm #ElectionNight
PinaSally|G_Eazy|0.7644|0.0|0.752|0.248|"RT @G_Eazy: PLEASE GO OUT AND VOTE WHATEVER YOU DO, THIS COULD BE THE MOST IMPORTANT ELECTION OF OUR LIVES #imwithher #fuckdonaldtrump"
HENRYFOREROJ|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
HENRYFOREROJ|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
Kilopher|IZOD|0.296|0.0|0.885|0.115|RT @IZOD: Share your voice this election. Make a statement with #MyVote2016 and Ken Bone in a red sweater. https://t.co/QX9fLqDpAL
Kilopher|twitter|0.296|0.0|0.885|0.115|RT @IZOD: Share your voice this election. Make a statement with #MyVote2016 and Ken Bone in a red sweater. https://t.co/QX9fLqDpAL
TransAmTobi|suttonimpaQt|0.3612|0.0|0.828|0.172|RT @suttonimpaQt: This election is like going outside to pick ya own switch.
ELau_87|THR|0.6369|0.0|0.625|0.375|RT @THR: Hollywood's best #Election2016 tweets https://t.co/FJx6s6ouYO https://t.co/PmPwzeyzE4
ELau_87|hollywoodreporter|0.6369|0.0|0.625|0.375|RT @THR: Hollywood's best #Election2016 tweets https://t.co/FJx6s6ouYO https://t.co/PmPwzeyzE4
MattZelinsky|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
MattZelinsky|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
kmrapp_7|Anna_Brodnik|0.0772|0.0|0.885|0.115|RT @Anna_Brodnik: I just want everyone to shut up about this election
LottNctc|chroniclelive|0.0|0.0|1.0|0.0|US presidential election: Results from New York - primary school North Tyneside  https://t.co/0fA9whgheA
deplorabletexas|OnlineMagazin|-0.5859|0.192|0.808|0.0|RT @OnlineMagazin:  #USA: Election Fraud by George #Soros-owned voting machine on Election Day in #Pennsylvania. #usaelections2016 #Sor
jgscroggins||0.0|0.0|1.0|0.0|"Your election PSA: sign up @ https://t.co/vxL0ZxUudQ. They will text or email you, or both, any time an election is in your area. #TurboVote"
jgscroggins|turbovote|0.0|0.0|1.0|0.0|"Your election PSA: sign up @ https://t.co/vxL0ZxUudQ. They will text or email you, or both, any time an election is in your area. #TurboVote"
bearoserod|BuzzFeedNews|-0.7028|0.271|0.729|0.0|"RT @BuzzFeedNews: 29 Most WTF Moments Of The Election: Hillary's Trump ""Joke"" #ElectionDay https://t.co/PNF7xkBxgB"
bearoserod|twitter|-0.7028|0.271|0.729|0.0|"RT @BuzzFeedNews: 29 Most WTF Moments Of The Election: Hillary's Trump ""Joke"" #ElectionDay https://t.co/PNF7xkBxgB"
LeLienDT|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
LeLienDT|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
biabru09|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
WilliamAmos|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
WilliamAmos|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
newsbreak|cnn|0.0|0.0|1.0|0.0|#cnn #Pantsuitnation goes to the polls: Women across the nation are wearing pantsuits on https://t.co/22fMeypy8W
havoksdemon|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
havoksdemon|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
garbagepanda|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
KneesaTata|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
Betweenthehedge|benshapiro|0.0|0.0|1.0|0.0|"RT @benshapiro: Our live coverage begins momentarily here -- with @andrewklavan, Jeremy Boreing, and a cast of thousands! https://t.co/l8gU"
Betweenthehedge|t|0.0|0.0|1.0|0.0|"RT @benshapiro: Our live coverage begins momentarily here -- with @andrewklavan, Jeremy Boreing, and a cast of thousands! https://t.co/l8gU"
xBenJamminx|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
CrumWillum|twitter|0.6166|0.0|0.598|0.402|Here is my election night....    :D https://t.co/lHFl0nYqND
remembermeoz|damianmcginty|0.4201|0.0|0.782|0.218|RT @damianmcginty: I am absolutely ready for this election to be over.
garth_wickham|SidneyCrosbyEgo|0.765|0.0|0.752|0.248|RT @SidneyCrosbyEgo: The best part about election day is that we get to watch McDavid and Crosby play before the world ends.
RyanWoodDFW|wusa9!|0.0|0.0|1.0|0.0|Election night at @wusa9!  @joanievas and I are heading up central coverage for @TEGNA!   https://t.co/xRLd5ymMxl
RyanWoodDFW|twitter|0.0|0.0|1.0|0.0|Election night at @wusa9!  @joanievas and I are heading up central coverage for @TEGNA!   https://t.co/xRLd5ymMxl
PublicBFLO|PublicBFLO|0.0|0.0|1.0|0.0|Tonight @PublicBFLO columnist Bruce Fisher will be doing election analysis on @WKBW. Tune in at 7:30! #ElectionNight
RF_Fayad|HuffPostPol|0.4215|0.147|0.58|0.272|RT @HuffPostPol: This election was colossally dumb and we're all lucky we survived it https://t.co/xFLKuRqNmn https://t.co/OiHLgURoiC
RF_Fayad|m|0.4215|0.147|0.58|0.272|RT @HuffPostPol: This election was colossally dumb and we're all lucky we survived it https://t.co/xFLKuRqNmn https://t.co/OiHLgURoiC
scottsaxton|Justin__West|0.0|0.0|1.0|0.0|"@Justin__West @AshleaOnAir Isn't it election ""afternoon"" for you?"
piwakawakaracin|TheSpinoffTV|0.0|0.0|1.0|0.0|"RT @TheSpinoffTV: The Spinoff Expert Panel will be updating every few seconds with the latest results, projections &amp; what have you.https:/"
jkoskenkorva|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
PatrickMillsaps|benparr|0.0|0.0|1.0|0.0|RT @benparr: How bots influenced the 2016 election: https://t.co/ncFcSeOMW5
PatrickMillsaps|refinery29|0.0|0.0|1.0|0.0|RT @benparr: How bots influenced the 2016 election: https://t.co/ncFcSeOMW5
Dreamy_Eyes5|twitter|0.6369|0.0|0.656|0.344|Best tweet I've seen about the election yet https://t.co/BWXmkL5ngI
JimmyBramlett|bpmoritz|0.0|0.0|1.0|0.0|RT @bpmoritz: Pizza is filtering into newsrooms around the country. Eyes are rolling in adjacent sports departments. https://t.co/60ORNPGmfy
JimmyBramlett|sportsmediaguy|0.0|0.0|1.0|0.0|RT @bpmoritz: Pizza is filtering into newsrooms around the country. Eyes are rolling in adjacent sports departments. https://t.co/60ORNPGmfy
TyBatiste|PittsburghPG|0.0|0.0|1.0|0.0|RT @PittsburghPG: Stay tuned to the Post-Gazette tonight for live local and national election results #pgvote2016 https://t.co/EKNIeOgPSZ h
TyBatiste|newsinteractive|0.0|0.0|1.0|0.0|RT @PittsburghPG: Stay tuned to the Post-Gazette tonight for live local and national election results #pgvote2016 https://t.co/EKNIeOgPSZ h
felipian|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
felipian|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
Jonnyboy_6969|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
buckitman|michaelharrisdr|0.4404|0.0|0.805|0.195|"RT @michaelharrisdr: #TrumpWinsBecause  says Patriots' Tom #Brady, Bill #Belichick supporting him @CNNPolitics https://t.co/kCFsGmSkPc"
buckitman|edition|0.4404|0.0|0.805|0.195|"RT @michaelharrisdr: #TrumpWinsBecause  says Patriots' Tom #Brady, Bill #Belichick supporting him @CNNPolitics https://t.co/kCFsGmSkPc"
kanjiklubs|Iitcompanys|-0.3265|0.142|0.761|0.096|RT @Iitcompanys: this election is so scary like some of y'all don't realize that almost everything that happens in the US affects the rest
cxrlittx|CNN|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
cxrlittx|twitter|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
_marhar|aislingd1989|0.743|0.0|0.769|0.231|@aislingd1989 Samantha Bee's coverage of the election has been A*. I'm aiming for 4am unless it's clear hilz has already won by then 
erickaa_zz|lizakoshyisbabe|-0.4404|0.266|0.734|0.0|RT @lizakoshyisbabe: Is anyone else scared about this election?
JamesWynn14|HRC4Prison|-0.296|0.136|0.864|0.0|RT @HRC4Prison: But Obama said there's no such thing as election fraudhttps://t.co/f7lP48RGlm #Wikileaks #PodestaEmails #ElectionFraud
sydawei|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
feministlawprof|twitter|0.0|0.0|1.0|0.0|"Getting this PowerPoint for tomorrow's Gender and Society class done before election results start rolling in, beca https://t.co/WDAv6vSEcq"
Humdingerding|NRO|0.0|0.0|1.0|0.0|"RT @NRO: Early Exit Polls: Trump Opens YUGE Gap between College-Educated, Non-College-Educated Whiteshttps://t.co/ADpCNhYfiC #ElectionNight"
vekmar|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
barjoriemerman|brokeymcpoverty|0.6705|0.0|0.593|0.407|thank goodness for @brokeymcpoverty leading me through this election night 
littledominguez|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
Momma__Kush|realDonaldTrump|0.4588|0.112|0.647|0.241|The thought of that trash @realDonaldTrump winning tonight is literally making my stomach upset. This election is a joke.
SixThreeOneFive|AriaWilsonGOP|-0.6884|0.226|0.774|0.0|RT @AriaWilsonGOP: Florida Election Worker Went Public With Massive Voter Fraud GOING DOWN RIGHT NOW!!! https://t.co/o1xK4N76gP https://t.c
SixThreeOneFive|everynewshere|-0.6884|0.226|0.774|0.0|RT @AriaWilsonGOP: Florida Election Worker Went Public With Massive Voter Fraud GOING DOWN RIGHT NOW!!! https://t.co/o1xK4N76gP https://t.c
AStageShout|GinnyMcQueen|-0.34|0.107|0.893|0.0|"RT @GinnyMcQueen: It's crazy to think that 2016 is our first election without a white, male candidate. What a time to be alive.#ImWithHer"
DireHeartbeat|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
grayy_ayshia|susanacaito19|-0.4101|0.199|0.801|0.0|RT @susanacaito19: this election is making me so nervous that I'm nauseous
laurenkierra|Lundentownn_|-0.2501|0.161|0.75|0.089|RT @Lundentownn_: Checking in on the election is like checking my bank account after a night out. I really don't want to see it and dread t
jensbachem|bbc|-0.4404|0.182|0.818|0.0|"Jeez... Once a fool, always a... ""George W Bush 'voted for none of the above'"" https://t.co/BSaKSLpOPy."
JustGoForIt|skyhookmike|-0.7254|0.272|0.728|0.0|RT @skyhookmike:  Because no REAL man WANTED that FILTHY MOUTH on their DI#%! Madonna Won't Honor Promise to Fellate Hillary Voter https:/
JustGoForIt||-0.7254|0.272|0.728|0.0|RT @skyhookmike:  Because no REAL man WANTED that FILTHY MOUTH on their DI#%! Madonna Won't Honor Promise to Fellate Hillary Voter https:/
CPCB|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
CPCB|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
_cpatrice|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
_cpatrice|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
BIGMONEYMETTA|UpshotNYT|0.5859|0.0|0.725|0.275|RT @UpshotNYT: When will we know we have a winner? https://t.co/1pMJXK7mS4 https://t.co/B87hwbBQZy
BIGMONEYMETTA|nytimes|0.5859|0.0|0.725|0.275|RT @UpshotNYT: When will we know we have a winner? https://t.co/1pMJXK7mS4 https://t.co/B87hwbBQZy
fergesor|hrtablaze|0.9207|0.0|0.645|0.355|RT @hrtablaze: My Bernie Sanders loving nephew who has been messing with me all election just told me he voted TRUMP !!! WOOT WOOT ! #elect
alyrose|jessicaseaman|0.0|0.0|1.0|0.0|RT @jessicaseaman: In the newsroom we have pizza for election night along with some cheese  dip   @alyrose https://t.co/Rq25rRo7zU
alyrose|twitter|0.0|0.0|1.0|0.0|RT @jessicaseaman: In the newsroom we have pizza for election night along with some cheese  dip   @alyrose https://t.co/Rq25rRo7zU
bleudawn7|alicebonasio|-0.5423|0.2|0.8|0.0|RT @alicebonasio: Millennials: get off your ass and #VOTEHILLARY NOW https://t.co/VlfdwzM0LX  #ElectionFinalThoughts #Election2016 @qz #br
bleudawn7|qz|-0.5423|0.2|0.8|0.0|RT @alicebonasio: Millennials: get off your ass and #VOTEHILLARY NOW https://t.co/VlfdwzM0LX  #ElectionFinalThoughts #Election2016 @qz #br
ThePhoenixFlare|julia_bergeron|0.6705|0.0|0.686|0.314|RT @julia_bergeron: Please let tonights election day sunset usher in a peaceful night. @SpaceCoastSkies https://t.co/wwOqRh0zpg
ThePhoenixFlare|twitter|0.6705|0.0|0.686|0.314|RT @julia_bergeron: Please let tonights election day sunset usher in a peaceful night. @SpaceCoastSkies https://t.co/wwOqRh0zpg
bellasmile2|CNET|0.0|0.0|1.0|0.0|RT @CNET: 5 live streams to watch if you're burnt out on the election #ElectionDay https://t.co/4Nk1jfeiHb
bellasmile2|twitter|0.0|0.0|1.0|0.0|RT @CNET: 5 live streams to watch if you're burnt out on the election #ElectionDay https://t.co/4Nk1jfeiHb
JarrodSHagenman|Variety|-0.8176|0.362|0.638|0.0|@Variety assholes.  That's automatic vote for Trump. Leave it to three #bushes to fuck up an election #imwithher
nwjerseyliz|CNN|0.4019|0.0|0.863|0.137|RT @CNN: Women across the nation are wearing pantsuits on #ElectionDay in support of Hillary Clinton https://t.co/TN3TeGDuDi #Pantsuitnatio
nwjerseyliz|cnn|0.4019|0.0|0.863|0.137|RT @CNN: Women across the nation are wearing pantsuits on #ElectionDay in support of Hillary Clinton https://t.co/TN3TeGDuDi #Pantsuitnatio
Tristan_runs|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
followtheAG|RealJamesWoods|0.0|0.0|1.0|0.0|RT @RealJamesWoods: This election in a nutshell... #Democrat #VoterFraud https://t.co/wFdlxex6UZ
followtheAG|twitter|0.0|0.0|1.0|0.0|RT @RealJamesWoods: This election in a nutshell... #Democrat #VoterFraud https://t.co/wFdlxex6UZ
murgaloo|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
meganvcolvin|JoshMarvine|0.7227|0.0|0.781|0.219|"RT @JoshMarvine: ""The iPhone doesn't have a headphone jack but the Galaxy literally explodes"" is a perfect metaphor for this election."
Laur_npr|samsanders|0.0|0.0|1.0|0.0|RT @samsanders: Here's @NPR's live election  night blog: https://t.co/UaPBLn1Kmu
Laur_npr|npr|0.0|0.0|1.0|0.0|RT @samsanders: Here's @NPR's live election  night blog: https://t.co/UaPBLn1Kmu
TheWillerix|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
deb_schiel|ABC|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
deb_schiel|abcnews|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
KevinMckechnie|RT_America|-0.4019|0.153|0.847|0.0|"RT @RT_America: BREAKING: Polling station on lockdown after shooting leaves 2 injured in Azuza, CA https://t.co/G0cuZ0bfH0 https://t.co/ffi"
KevinMckechnie|rt|-0.4019|0.153|0.847|0.0|"RT @RT_America: BREAKING: Polling station on lockdown after shooting leaves 2 injured in Azuza, CA https://t.co/G0cuZ0bfH0 https://t.co/ffi"
ohcrapstyles|HSupdating|0.5948|0.0|0.819|0.181|"RT @HSupdating: In honor of Election Day in America, never forget when Harry was rumored to be having an affair with Barack Obama. https://"
ohcrapstyles||0.5948|0.0|0.819|0.181|"RT @HSupdating: In honor of Election Day in America, never forget when Harry was rumored to be having an affair with Barack Obama. https://"
jefecich|twitter|0.0|0.0|1.0|0.0|Election Day #FoxNews2016 #ElectionNight #Vote2016 #NBC2016 https://t.co/jlUrnFCdJD
mckbrowny|OllyNewport|0.4019|0.0|0.787|0.213|RT @OllyNewport: Just preparing for my election party tonight. #Election2016 https://t.co/8b2SVmbmTZ
mckbrowny|twitter|0.4019|0.0|0.787|0.213|RT @OllyNewport: Just preparing for my election party tonight. #Election2016 https://t.co/8b2SVmbmTZ
PvillePostNews|weebly|0.0|0.0|1.0|0.0|Check out our newest blog post! #electionnight #democrats #republicans https://t.co/1mD2uGMOJa via @weebly
PvillePostNews|thepleasantvillepost|0.0|0.0|1.0|0.0|Check out our newest blog post! #electionnight #democrats #republicans https://t.co/1mD2uGMOJa via @weebly
mariaeke|bipartisanreport|0.2103|0.0|0.857|0.143|BREAKING: FBI STUNS America With Election Day Trump/Russia Warrant Announcement (DETAILS) https://t.co/MSmf7cvINR
OfficialYoungRB|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
OfficialYoungRB|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
CraigJ_NandO|twitter|0.4019|0.0|0.847|0.153|"We're all just hangin' out at the McCroy election night party, not yet underway. #ncpol https://t.co/LbrGlMYc8X"
lp_1516|El_Ma3stro77|0.0775|0.076|0.799|0.125|RT @El_Ma3stro77: @lp_1516 @IZOD I didn't vote you know that lol cause I know it's important to do it but I don't think it's worth in this
baygui|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
baygui|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
shar_veshh|BazK10|0.5719|0.0|0.73|0.27|RT @BazK10: I will eat this if trump wins the election  https://t.co/SGLHSg7MmO
shar_veshh|twitter|0.5719|0.0|0.73|0.27|RT @BazK10: I will eat this if trump wins the election  https://t.co/SGLHSg7MmO
into_thev0id|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
into_thev0id|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
Happy_Dais|BarnabyEdwards|0.5859|0.051|0.725|0.225|RT @BarnabyEdwards: It's hard to know who I'd vote for in the US election: the candidate backed by everyone I respect or the one endorsed b
kabbath|KHQA|0.0|0.0|1.0|0.0|RT @KHQA: Eric Trump illegally posts pic of completed NY ballot on Twitterhttps://t.co/o3ic19ZzeU
electricpac|mike_pence|0.0|0.0|1.0|0.0|"RT @mike_pence: This Election Day, America is standing at the crossroads of history. RT this if you're voting for @realDonaldTrump. Togethe"
LuckymeEva|BBCBreaking|0.9041|0.0|0.617|0.383|"RT @BBCBreaking: ""I'll do the very best I can if I'm fortunate enough to win today"" - @HillaryClinton casts her ballot #Election2016 https:"
ellie_gretter|parker_maurer|0.0|0.0|1.0|0.0|RT @parker_maurer: One of my biggest pet peeves throughout this election is how people are so quick to judge/bash someone based on who they
LeahVossVisuals|twitter|0.7959|0.0|0.664|0.336|The Noveaux Honkies are playing a free show until 8 p.m. at Terra Fermata at Crystal Lucas' election night party! https://t.co/19XtTXwzxv
fumiplagg|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Its Election Day and polls are officially open. When will you vote today? Confirm where to go here: https://t.co/jfd3C
fumiplagg|t|0.0|0.0|1.0|0.0|RT @HillaryClinton: Its Election Day and polls are officially open. When will you vote today? Confirm where to go here: https://t.co/jfd3C
CodeRedSME|instagram|0.0|0.0|1.0|0.0|"While waiting for the results of the election, eating cookies and drinking gin. #lenny&amp;larry's https://t.co/jRpqwZ8USI"
CollaurJohn|TheCanarySays|-0.0516|0.105|0.798|0.097|"RT @TheCanarySays: While all are fixated on the US election, an appalling truth about the UK has quietly been revealed https://t.co/cWI4o8S"
CollaurJohn|t|-0.0516|0.105|0.798|0.097|"RT @TheCanarySays: While all are fixated on the US election, an appalling truth about the UK has quietly been revealed https://t.co/cWI4o8S"
FehlJohn|TheLastRefuge2|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
FehlJohn|twitter|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
rivjudes|Maddynx|0.0|0.0|1.0|0.0|RT @Maddynx: Twitter on Election Dayhttps://t.co/04p0nkjyiw
Jonfromncl|mrchrisaddison|-0.4118|0.116|0.884|0.0|"RT @mrchrisaddison: The last time I was watching a US election this tense, I was standing in the room with Selina Meyer and her team."
ClockworkJest|tomlucy|0.6768|0.0|0.791|0.209|RT @tomlucy: I'm excited about the US election but it's the sort of excitement you get before you put a knife in the toaster.
AndreHeadlee|nytimes|0.0|0.0|1.0|0.0|Presidential Election Results https://t.co/hBDPoYigk0
PTLHayward|clydesdalequeen|0.0|0.0|1.0|0.0|RT @clydesdalequeen: Feel for my USA teacher peeps..rationalizing this election with kids. May have an ulcer b/f it's over and I'm Cdn ! #
varunpramanik|JonErlichman|0.0|0.0|1.0|0.0|RT @JonErlichman: Things that didn't exist election night in 2008:UberiPadInstagramSnapchatWhatsAppPinterestPeriscopeOculusSlack
geek4fun|veggienut|-0.2732|0.163|0.724|0.113|RT @veggienut: Dog took a shit in the living room so now I think I'm ready for Election coverage. https://t.co/DGMEv1eop1
geek4fun|twitter|-0.2732|0.163|0.724|0.113|RT @veggienut: Dog took a shit in the living room so now I think I'm ready for Election coverage. https://t.co/DGMEv1eop1
patriciayingst|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
patriciayingst|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
canderson1989|girlsreallyrule|0.3612|0.0|0.839|0.161|@girlsreallyrule Election night event in NYC. Ready to shatter the glass. #ElectionNight #ImWithHer https://t.co/QneFY90TDG
canderson1989|twitter|0.3612|0.0|0.839|0.161|@girlsreallyrule Election night event in NYC. Ready to shatter the glass. #ElectionNight #ImWithHer https://t.co/QneFY90TDG
JSara1234|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
seufert|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
seufert|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
MollyQuilitzsch|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
MollyQuilitzsch|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
ReneeLoder|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
ReneeLoder|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
nothing_exists|chrislhayes|-0.5256|0.159|0.841|0.0|RT @chrislhayes: Trump is already laying the groundwork to contest the legitimacy of the election and it's incredibly dangerous.
chipgw|ToryBelleci|0.0|0.0|1.0|0.0|RT @ToryBelleci: It's Election Night! Let the results pour in. #election2016 https://t.co/aaynBMS2uU
chipgw|instagram|0.0|0.0|1.0|0.0|RT @ToryBelleci: It's Election Night! Let the results pour in. #election2016 https://t.co/aaynBMS2uU
libsidcap|akcdogloversNeed|0.0|0.0|1.0|0.0|@akcdoglovers:Need break from election coverage?We've got just thing!https://t.co/fF0f6LIG1l #dogs #doglover #cute https://t.co/OvT6gTIDfc
libsidcap|akc|0.0|0.0|1.0|0.0|@akcdoglovers:Need break from election coverage?We've got just thing!https://t.co/fF0f6LIG1l #dogs #doglover #cute https://t.co/OvT6gTIDfc
CarlosIsCarLost|MaduroOfficial|0.0|0.0|1.0|0.0|RT @MaduroOfficial: USA ELECTION UPDATEDonald Trump -   22.4%Hilary Clinton -   16.6%PSUV.               -  61.1%
2camxxx|barnabybabybump|0.0|0.0|1.0|0.0|RT @barnabybabybump: got my election sticker for tomorrow https://t.co/QQ6myPejGO
2camxxx|twitter|0.0|0.0|1.0|0.0|RT @barnabybabybump: got my election sticker for tomorrow https://t.co/QQ6myPejGO
schafedog12|CharlieDayQuote|0.0|0.0|1.0|0.0|RT @CharlieDayQuote: After the election results tonight... https://t.co/cmPwW4Jded
schafedog12|twitter|0.0|0.0|1.0|0.0|RT @CharlieDayQuote: After the election results tonight... https://t.co/cmPwW4Jded
Grammy8|TeaPartyOrg|-0.5574|0.217|0.783|0.0|RT @TeaPartyOrg: 2 Florida Election Officials Fired For Not Adhering To Procedure And Policy - https://t.co/nrcxcYAy7y
Grammy8|teaparty|-0.5574|0.217|0.783|0.0|RT @TeaPartyOrg: 2 Florida Election Officials Fired For Not Adhering To Procedure And Policy - https://t.co/nrcxcYAy7y
jasonnellis|melissaFTW|0.128|0.0|0.914|0.086|RT @melissaFTW: We all deserve a Purge-like rule where the day after the election every drug is legal.
luletobe|SunSentinel|-0.4019|0.162|0.838|0.0|"RT @SunSentinel: Election 2016: Voters face machine problems, long lines in some states https://t.co/U3XvoCCPQj https://t.co/oMHXLsTv8o"
luletobe|sun-sentinel|-0.4019|0.162|0.838|0.0|"RT @SunSentinel: Election 2016: Voters face machine problems, long lines in some states https://t.co/U3XvoCCPQj https://t.co/oMHXLsTv8o"
ohhbrynn|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
ohhbrynn|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
HickmanJessie|breanna_owenss|-0.7358|0.342|0.658|0.0|RT @breanna_owenss: I WANNA SAY SO MANY BAD WORDS ABOUT THIS ELECTION 
TeamCrazyMatt|FiveThirtyEight|0.1027|0.115|0.752|0.133|RT @FiveThirtyEight: Preliminary exit polls show that many voters were motivated by dislike of one of the candidates. https://t.co/0soCpm3M
TeamCrazyMatt|t|0.1027|0.115|0.752|0.133|RT @FiveThirtyEight: Preliminary exit polls show that many voters were motivated by dislike of one of the candidates. https://t.co/0soCpm3M
lexi_havel97|MaggieBecka|0.0258|0.113|0.769|0.117|RT @MaggieBecka: i am freaking the heck out over this election. i cannot understand why anyone would think trump would be a good leader
tlynn561|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
tlynn561||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
Alexiaa_Minaj|FrankLuntz|0.4019|0.0|0.891|0.109|"RT @FrankLuntz: All eyes will be in Virginia for 2017.Tim Kaine's Senate seat will open up, and they will have a special election.  #Elec"
elostris|theguardian|0.0|0.0|1.0|0.0|us presidential elections 101 https://t.co/Azn03z7dC3
taytay007007007|HalleyBorderCol|0.7703|0.0|0.74|0.26|"RT @HalleyBorderCol: For anyone wanting election results as them come in, the Guardian site seems quite good. Looking good for #Trump!htt"
LouiseDoire|MiamiHerald|0.3818|0.0|0.852|0.148|"RT @MiamiHerald: On Election Day, the Miami Herald's Editorial Page makes a bold statement: ENOUGH SAID. https://t.co/RrUKzCgdDx"
LouiseDoire|twitter|0.3818|0.0|0.852|0.148|"RT @MiamiHerald: On Election Day, the Miami Herald's Editorial Page makes a bold statement: ENOUGH SAID. https://t.co/RrUKzCgdDx"
HometownHero81|MattMoretta|0.8934|0.0|0.545|0.455|"RT @MattMoretta: Plot twist: Matthew McConaughey wins election, everyone receives a brand new Lincoln, happiness is restored alright alrigh"
marthajadams|AAUW|-0.3595|0.122|0.878|0.0|RT @AAUW: THIS! These Black Women Also Deserve A Visit To Their Graves On Election Day: https://t.co/6N40THpHOr? #ElectionDay #ItsMyVote by
marthajadams|huffingtonpost|-0.3595|0.122|0.878|0.0|RT @AAUW: THIS! These Black Women Also Deserve A Visit To Their Graves On Election Day: https://t.co/6N40THpHOr? #ElectionDay #ItsMyVote by
webcentraltv|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
webcentraltv|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
elizabethfais|CatFoodBreath|0.6996|0.0|0.721|0.279|RT @CatFoodBreath: Looks like a 4-way race in the election for favorite CFB character! #Vote2016 22%Thing Two25%Nativity Sheep28%Labradu
gollottomarco|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
gollottomarco|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
numinouscosmos|youtube|0.0|0.0|1.0|0.0|2016 ELECTION PLAYLIST - USSR NATIONAL ANTHEM:https://t.co/5aHE98yQFA
Roryyy_b|bet365|0.8225|0.0|0.703|0.297|Get trump to win the election at 9/2 or Clinton 1/6Underdog got the brexit win will it happen again? https://t.co/zvD2gTWU4I
mijsetay|truthout|0.4939|0.0|0.814|0.186|RT @truthout: Today's Election Results Could Affect Mental Health Care for Millions https://t.co/m0po3UGBAT #ElectionDay #mentalhealth
mijsetay|truth-out|0.4939|0.0|0.814|0.186|RT @truthout: Today's Election Results Could Affect Mental Health Care for Millions https://t.co/m0po3UGBAT #ElectionDay #mentalhealth
Str8Grandmother|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
Str8Grandmother||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
helenjowens|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
TheJLoSpot|twitter|-0.8856|0.378|0.537|0.085|I'm glad the judge stopped this fat ugly racist orange oompa loompa piece of shit!! He'd only use it to lie &amp; say t https://t.co/c85xCTipJe
ukiparmy|WDFx2EU8|-0.1531|0.121|0.781|0.098|"RT @WDFx2EU8: The  election in a nutshell. On the left, Lady Gaga dancing like a dipshit at Clinton concert. On right, Mike Pence talking a"
elliegallgher21|Things4WhitePpl|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
elliegallgher21|twitter|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
MrMcGov|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
MrMcGov|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
VoteTrumpPence7|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
donna_heinrich|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
Guille_Roma|lord_iniesta|0.0|0.0|1.0|0.0|@lord_iniesta https://t.co/NdTJud6mz4 real time
Guille_Roma|politico|0.0|0.0|1.0|0.0|@lord_iniesta https://t.co/NdTJud6mz4 real time
mal_FUNK_tion|briankoppelman|0.3612|0.0|0.906|0.094|RT @briankoppelman: Karl Rove back on Fox News election night after the debacle 4 yrs ago would be like me sitting down to write Runner Run
davo_iguodala|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
davo_iguodala|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
CKlein5852|AdamsFlaFan|-0.128|0.215|0.633|0.152|RT @AdamsFlaFan: Hero Judge Stands Up For Democracy And Rejects Trump's Nevada Election Day Lawsuit via @politicususa https://t.co/v32RI9gi
CKlein5852|t|-0.128|0.215|0.633|0.152|RT @AdamsFlaFan: Hero Judge Stands Up For Democracy And Rejects Trump's Nevada Election Day Lawsuit via @politicususa https://t.co/v32RI9gi
NickKlopsis|Newsday|0.0|0.0|1.0|0.0|"While some people wait in line to vote, @Newsday waits in line for election night subs. https://t.co/8ulNTJqtU4"
NickKlopsis|twitter|0.0|0.0|1.0|0.0|"While some people wait in line to vote, @Newsday waits in line for election night subs. https://t.co/8ulNTJqtU4"
MikeConnors|SheenaGoodyear|0.3612|0.0|0.828|0.172|RT @SheenaGoodyear: Not working on election night makes me feel like such a muggle.
gaelicdiana|michaelbeatty3|0.0|0.0|1.0|0.0|RT @michaelbeatty3: If you're whipping out the Khan family on election night...You are scared....#electionday #MAGA https://t.co/0J68VGtm
gaelicdiana|t|0.0|0.0|1.0|0.0|RT @michaelbeatty3: If you're whipping out the Khan family on election night...You are scared....#electionday #MAGA https://t.co/0J68VGtm
kirsmu|JinkxMonsoon|0.9392|0.0|0.578|0.422|"RT @JinkxMonsoon: Here I am the first time Obama won, with my friend Samie doing enough celebrating for the two of us! Happy Election Day e"
rbxlifestyle|KathleenLights1|0.4199|0.141|0.573|0.286|RT @KathleenLights1: Hope everyone voted today! This election has traumatized me.... I pray for America.
Alyssa_trapani|jesssmauro|-0.6369|0.174|0.826|0.0|RT @jesssmauro: This election has made so many people turn against each other. People are becoming divided and filled with hatred
dggabber|ilnews|0.0|0.0|1.0|0.0|Election day in Illinois: What's at stake? - Illinois News Network https://t.co/uvMsV05E47
agent_it|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
agent_it|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
rkellett|twitter|0.6249|0.0|0.709|0.291|What it takes to make it great on election night https://t.co/FZu5sf2Dcc
RMarcelc|wesearchr|0.6633|0.0|0.811|0.189|"RT @wesearchr: To collect our $6720 REWARD for documented proof of #ElectionFraud, SUBMIT IT to the page here: https://t.co/ThS6MrnNCF #MAG"
RMarcelc|wesearchr|0.6633|0.0|0.811|0.189|"RT @wesearchr: To collect our $6720 REWARD for documented proof of #ElectionFraud, SUBMIT IT to the page here: https://t.co/ThS6MrnNCF #MAG"
thewhiteflame21|ESPNStatsInfo|0.34|0.0|0.906|0.094|RT @ESPNStatsInfo: Connor McDavid &amp; Sidney Crosby meet for 1st timeMario Lemieux &amp; Wayne Gretzky played vs each other for 1st time on Ele
RickOsborne2|WordSmithGuy|0.0|0.0|1.0|0.0|RT @WordSmithGuy: Florida Panhandle &amp; Michigan: You have 1 hour &amp; 15 minutes to make history. This entire election may be decided by you gu
twt6969|globeandmail|0.0772|0.0|0.949|0.051|"RT @globeandmail: #ElectionDay is going to be a long one. If all you want to know is when the results will be announced, here you gohttps:"
fatimaaCakess|biggabossben|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
fatimaaCakess|twitter|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
ch1election|WSBT|-0.4019|0.213|0.787|0.0|RT @WSBT: Live video from battleground state of New Hampshire: https://t.co/JUgiX5tUYP
ch1election|wsbt|-0.4019|0.213|0.787|0.0|RT @WSBT: Live video from battleground state of New Hampshire: https://t.co/JUgiX5tUYP
EfrataAxayaRosa|ReutersTV|0.0|0.0|1.0|0.0|RT @ReutersTV: #Election2016: The trail and the tumult https://t.co/mmpNiISEp4 https://t.co/yQZXwqCBV5
EfrataAxayaRosa|app|0.0|0.0|1.0|0.0|RT @ReutersTV: #Election2016: The trail and the tumult https://t.co/mmpNiISEp4 https://t.co/yQZXwqCBV5
scelzi_dolores|StacyBrewer18|0.0|0.0|1.0|0.0|RT @StacyBrewer18: 2016 Election Day: Live Updates - Breitbart https://t.co/ppsyYS9fdP
scelzi_dolores|linkis|0.0|0.0|1.0|0.0|RT @StacyBrewer18: 2016 Election Day: Live Updates - Breitbart https://t.co/ppsyYS9fdP
NickDawybida|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
loveloso_|DarkerThanAkon|0.0|0.0|1.0|0.0|RT @DarkerThanAkon: IT'S ELECTION DAY I KNOW YA'LL WILL MAKE THE RIGHT DECISION https://t.co/yF73IzfIk4
loveloso_|twitter|0.0|0.0|1.0|0.0|RT @DarkerThanAkon: IT'S ELECTION DAY I KNOW YA'LL WILL MAKE THE RIGHT DECISION https://t.co/yF73IzfIk4
hckysnyder|oliviarlaborde|0.8346|0.0|0.583|0.417|RT @oliviarlaborde: hey @realDonaldTrump u better win so I can vote for u next election!!!!!!! @sgmauldin
magicisalways|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
magicisalways|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Yonna_Ziel|lesleythornton_|-0.7939|0.252|0.748|0.0|RT @lesleythornton_: its really disgusting and sad the way some people minds work ... and it all came out during this presidential election
Beerad30|TheSeigeDFS|0.7096|0.0|0.734|0.266|"RT @TheSeigeDFS: Hope this election is the final straw America needs to remember that primaries matter, we should have better options than"
Kbabyymota|TeaBaggett|0.4019|0.0|0.87|0.13|"RT @TeaBaggett: After this election I will be hosting an ""End of the World"" party. Rt if you wanna come"
JoshAmos96|Amy_ninetyeight|0.5574|0.0|0.69|0.31|@Amy_ninetyeight Nothing beats his general election swing ones hahaha
KWebb_Harward|__Weston__|0.2263|0.193|0.541|0.266|"RT @__Weston__: The world fails to realize that no matter who wins the election, God will remain in control."
IOM_USA|H_NAILI|0.0|0.0|1.0|0.0|RT @H_NAILI: Tonight 1st Muslim refugee &amp; 1st Somali American woman to hold elected office in US could be elected https://t.co/bONTI2WyuA #
IOM_USA|theguardian|0.0|0.0|1.0|0.0|RT @H_NAILI: Tonight 1st Muslim refugee &amp; 1st Somali American woman to hold elected office in US could be elected https://t.co/bONTI2WyuA #
mazzy0108|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
mazzy0108|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
hunter_ripley|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
SoyerJanis|athena_Insight|0.0|0.0|1.0|0.0|RT @athena_Insight: Medical marijuana is on the ballot in #Florida. See how it may affect #opioid prescribing rates. #election https://t.co
SoyerJanis|t|0.0|0.0|1.0|0.0|RT @athena_Insight: Medical marijuana is on the ballot in #Florida. See how it may affect #opioid prescribing rates. #election https://t.co
notericisboss84|BoofBaldy|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
notericisboss84|twitter|0.5859|0.0|0.774|0.226|"RT @BoofBaldy: ""And the winner of the 2016 presidential election is... Donald Trump""Immigrants: https://t.co/kpC1BvnFSL"
cchsctv|facebook|0.0|0.0|1.0|0.0|CTV Teens Vote 7PMCTV Election Coverage https://t.co/Nqn5midjrg
Hanto38Le|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
Hanto38Le|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
KristinaF1977|FreddieCampion|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
KristinaF1977|twitter|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
CarusiPrincipal|CarusiMS|0.0258|0.0|0.939|0.061|RT @CarusiMS: 8th Grade Election Night tonight 7-9pm. Enter through Gym lobby and go to our cafeteria. https://t.co/biG7KAwcnm
CarusiPrincipal|twitter|0.0258|0.0|0.939|0.061|RT @CarusiMS: 8th Grade Election Night tonight 7-9pm. Enter through Gym lobby and go to our cafeteria. https://t.co/biG7KAwcnm
jkbriseno|nytimes|0.5859|0.0|0.725|0.275|RT @nytimes: When will we know when we have a winner? https://t.co/58YOEs664i
jkbriseno|nytimes|0.5859|0.0|0.725|0.275|RT @nytimes: When will we know when we have a winner? https://t.co/58YOEs664i
Aspennicole17|precious_oxox|-0.6169|0.314|0.686|0.0|RT @precious_oxox: this election is fucking with my anxiety. Donald Trump cannot win.
ramesh_tnt|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
ramesh_tnt|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
Axellent33|Verge|0.5106|0.0|0.708|0.292|Donald Trump's website enjoyed a brief democracy https://t.co/y7zBMbqU8i via @Verge
Axellent33|theverge|0.5106|0.0|0.708|0.292|Donald Trump's website enjoyed a brief democracy https://t.co/y7zBMbqU8i via @Verge
tzraik|WSJ|0.2023|0.0|0.917|0.083|"RT @WSJ: Election night guide: The top things to watch, with key times and races of the night https://t.co/l6LIuGSM0f #election2016  https"
tzraik|blogs|0.2023|0.0|0.917|0.083|"RT @WSJ: Election night guide: The top things to watch, with key times and races of the night https://t.co/l6LIuGSM0f #election2016  https"
AmyBlankenship|BenNadel|0.5473|0.0|0.665|0.335|@BenNadel Post-Election: Game of Thrones binge watch LOL
gregmroscoe|MayorOfLA|0.8478|0.0|0.674|0.326|"RT @MayorOfLA: The importance of this election is too great to simply stay home. Please get out and vote, LA! Visit https://t.co/277rgwAQLs"
gregmroscoe|lavote|0.8478|0.0|0.674|0.326|"RT @MayorOfLA: The importance of this election is too great to simply stay home. Please get out and vote, LA! Visit https://t.co/277rgwAQLs"
AlanbNYC|twitter|0.6105|0.108|0.505|0.387|Ok this is funny. A little humor I suspect is needed on election day  https://t.co/6F6O91hsZP
CDNutz14|Livestream|0.0|0.0|1.0|0.0|Watch Election 2016 Livestream on @Livestream: https://t.co/Ebsdg2TceU
CDNutz14|livestream|0.0|0.0|1.0|0.0|Watch Election 2016 Livestream on @Livestream: https://t.co/Ebsdg2TceU
mdavkes|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
mdavkes|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
HiTechWorldNews|route|0.0|0.0|1.0|0.0|How likely is it for someone to hack the US election? https://t.co/VPE8lSn6jH https://t.co/Oflf6pdSC1
citroncool|dril|0.0|0.0|1.0|0.0|RT @dril: if you ask me this election could end about 100 different ways:1) trump gets 0% of the vote2) trump gets 1% of the vote3) trum
BookHoundsBlog|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
mohermes2020|DocFaustine|0.0|0.0|1.0|0.0|"RT @DocFaustine: Three o'clock in the morning and still awake, following US election results https://t.co/5DyTzdU4XC"
mohermes2020|instagram|0.0|0.0|1.0|0.0|"RT @DocFaustine: Three o'clock in the morning and still awake, following US election results https://t.co/5DyTzdU4XC"
artofwar73|CNN|0.4753|0.0|0.781|0.219|Watching @CNN election results likes it's a football playoff game!  Where's the popcorn?
marveItrade|mashable|0.0|0.0|1.0|0.0|RT @mashable: Caught! Donald Trump was peeking at his wife's election ballot  #ElectionNight https://t.co/1CsOJNnkpo
marveItrade|twitter|0.0|0.0|1.0|0.0|RT @mashable: Caught! Donald Trump was peeking at his wife's election ballot  #ElectionNight https://t.co/1CsOJNnkpo
BrendanTN_|RCDefense|0.0|0.0|1.0|0.0|RT @RCDefense: Cyberwarfare Amidst the U.S. #Election | @BrendanTN_ @LowyInstitute #ElectionDay #ElectionNight #Election2016 https://t.co/3
BrendanTN_|twitter|0.0|0.0|1.0|0.0|RT @RCDefense: Cyberwarfare Amidst the U.S. #Election | @BrendanTN_ @LowyInstitute #ElectionDay #ElectionNight #Election2016 https://t.co/3
thefiddleflores|HillaryClinton|0.4019|0.0|0.863|0.137|@HillaryClinton @HFA @katyperry @HillaryForNY this election party is fucking bs. I waited 3hrs 4 tix &amp; 10hrs @javitscenter. Can't c nothing.
ShekYerbouti|twitter|0.1071|0.102|0.764|0.134|I would like to call the election but I can't find their number https://t.co/c8LK3HoDdT
franklapore|politico|-0.5859|0.348|0.652|0.0|Trump seizes on isolated glitches to fuel rigged election claims  https://t.co/AVEY0b9tPT
FLMENFORTRUMP|SonofLiberty357|0.4939|0.0|0.824|0.176|RT @SonofLiberty357: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/VpmqCeml3e
FLMENFORTRUMP|thegatewaypundit|0.4939|0.0|0.824|0.176|RT @SonofLiberty357: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/VpmqCeml3e
BULGEBULL|t|0.0|0.0|1.0|0.0|WATCH LIVE: 5 Streaming News Channels Covering Election Night 2016 https://t.co/48zkTcOeYYIf youre looking for https://t.co/bAnUclGknV
e_poll2016|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
e_poll2016|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
Stepto|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
schwiick|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
schwiick|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
NaisBtd|CBCAlerts|-0.8481|0.326|0.674|0.0|"RT @CBCAlerts: One dead in shooting in California, three injured near polling station. No indication so far that it is election-related: re"
tlvrp_russia|therussophile|-0.2732|0.195|0.667|0.138|#Moscow #SaintPetersburg Stanford University Confirms Democratic 2016 Election Fraud In Favor of Hillary Clinton https://t.co/9Ps7WcZp6q
thvideogamenews|asunnydisposish|-0.2263|0.076|0.924|0.0|"RT @asunnydisposish: As someone who can't vote today but will still be affected by the election results, I urge you to not throw away your"
neyotherock|TrailerJamShow|-0.3182|0.15|0.85|0.0|RT @TrailerJamShow: The election is causing loads of accidents on the highway  #TrailerJamShow https://t.co/p5UNoTWqDN
neyotherock|twitter|-0.3182|0.15|0.85|0.0|RT @TrailerJamShow: The election is causing loads of accidents on the highway  #TrailerJamShow https://t.co/p5UNoTWqDN
IrwanFelany|instagram|0.4215|0.0|0.641|0.359|United State Election 2016#kamiawani #usaelections2016 https://t.co/VA9MS52JBm
Owfield|NewsHour|0.0|0.0|1.0|0.0|"RT @NewsHour: Whether you've yet to vote or have already voted, let us know why you cast a ballot in this election. Tell us with #MyVotePBS"
janet_cutts|Reuters|0.0|0.0|1.0|0.0|RT @Reuters: Democrats hold slight edge in contest to control Senate https://t.co/OAR9uCsY1B https://t.co/VviwIv3AqY
janet_cutts|reuters|0.0|0.0|1.0|0.0|RT @Reuters: Democrats hold slight edge in contest to control Senate https://t.co/OAR9uCsY1B https://t.co/VviwIv3AqY
AvoDead|VenomsDevil|0.0|0.0|1.0|0.0|@VenomsDevil voting isn't strictly presidential in America. There is a host of propositions and local voting on Election Day
kinkyseoks|PJMedia_com|0.0|0.0|1.0|0.0|RT @PJMedia_com: Vote: What will you be drinking while watching election returns tonight?#ElectionNight #voted
Koxinga8|breitbart|0.5859|0.0|0.774|0.226|Frank Luntz: #Trump Could Win Michigan  Working-Class Turnout 'Much Higher than Expected' - Breitbart https://t.co/gIclIzCOzS
FamousPixs|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
FamousPixs|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
TRUMPNEXTPRES16|RealBenCarson|0.5423|0.0|0.791|0.209|RT @RealBenCarson: Tomorrow's election is 'The Political Class' vs 'We The People.' Please read and share my newest article.https://t.co/
davedbody|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
davedbody|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
patriciayingst|WSJPolitics|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
patriciayingst|wsj|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
lillayyyy_|LKiddy2|0.0|0.0|1.0|0.0|RT @LKiddy2: If our founding fathers could see this election they'd probably give our country back to the British.
laceylfischer_|SoDamnTrue|0.3612|0.0|0.828|0.172|RT @SoDamnTrue: what twitter will be like today since its election day https://t.co/kVb11TM7CJ
laceylfischer_|vine|0.3612|0.0|0.828|0.172|RT @SoDamnTrue: what twitter will be like today since its election day https://t.co/kVb11TM7CJ
JOHNTFALVEYSR|RT_America|-0.7717|0.34|0.66|0.0|"RT @RT_America: BREAKING: Reports of one dead after gunman opened fire in Azusa, CA https://t.co/G0cuZ0bfH0"
JOHNTFALVEYSR|rt|-0.7717|0.34|0.66|0.0|"RT @RT_America: BREAKING: Reports of one dead after gunman opened fire in Azusa, CA https://t.co/G0cuZ0bfH0"
XaviVenegas|IZOD|0.296|0.0|0.833|0.167|RT @IZOD: America votes. Join the Election Day conversation with #MyVote2016 https://t.co/BWuiwAxas6
XaviVenegas|twitter|0.296|0.0|0.833|0.167|RT @IZOD: America votes. Join the Election Day conversation with #MyVote2016 https://t.co/BWuiwAxas6
karmunyu|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
karmunyu|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
grandmaKim27|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
Cyber_Legendary|twitter|0.3612|0.0|0.8|0.2|I'm ready for the results of the election. #electionday #ElectionNight https://t.co/iHMRf5yZcQ
tobibeth1|TheAnonnMessage|0.4003|0.0|0.77|0.23|@TheAnonnMessage Not determined if shooting is related to election yet!
TedFlintKansas|ericmichel|0.3612|0.0|0.857|0.143|RT @ericmichel: I am going to hate-watch CNN's election night coverage like the last season of Dexter
BULGEBULL|i2|0.4019|0.0|0.838|0.162|WATCH LIVE: Hillary Clinton and Donald Trump Hold Election Night Parties Only A Mile Apart  https://t.co/vGY5zOkGg6
curraheave|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
curraheave|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
Toastiewiththe|nytimes|0.5859|0.0|0.725|0.275|RT @nytimes: When will we know when we have a winner? https://t.co/58YOEs664i
Toastiewiththe|nytimes|0.5859|0.0|0.725|0.275|RT @nytimes: When will we know when we have a winner? https://t.co/58YOEs664i
LabourNHSJAN|independent|0.296|0.0|0.885|0.115|Eric Trump illegally shares photo of him voting for his dad to be president | The Independent - www.independent. https://t.co/oee14c9qiI
OdellSZN|StephForMVP30|0.7955|0.0|0.718|0.282|RT @StephForMVP30: If Trump or Hillary wins the election I'm moving out the country! Goodbye America and hello United States!
mariachooch|iHumbleThots|0.3612|0.0|0.737|0.263|RT @iHumbleThots: Waiting on Election results like https://t.co/4elYh2O7Ic
mariachooch|twitter|0.3612|0.0|0.737|0.263|RT @iHumbleThots: Waiting on Election results like https://t.co/4elYh2O7Ic
VZoey101|Khanoisseur|0.765|0.0|0.752|0.248|RT @Khanoisseur: Easily the best use of a campaign plane this election season: Clinton team (with Jon Bon Jovi) pull off a spectacular mann
PANKsinatra|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
PANKsinatra|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
hkmeehan|WDFx2EU8|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
hkmeehan|conservativeeagles|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
TheSpencerSapp|twitter|0.0|0.0|1.0|0.0|The only way I'll be able to get through the waning hours of the election... https://t.co/xJgPLv0FS9
laurie6805|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
laurie6805|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
hueDothanh|YouTube|0.0|0.0|1.0|0.0|Election 2016 Voting under way for next president: https://t.co/tUEDCcpImG qua @YouTube
hueDothanh|youtube|0.0|0.0|1.0|0.0|Election 2016 Voting under way for next president: https://t.co/tUEDCcpImG qua @YouTube
charissemarie|inquisitr|0.0|0.0|1.0|0.0|Get Live #Election Results Streaming Online And Be The First To Know Who The #President Is https://t.co/eDTWkHqQNF
zoomollogist|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
KweschnMedia|ajplus|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
KweschnMedia|twitter|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
dlmassepuh|RitaCosby|0.5374|0.0|0.852|0.148|RT @RitaCosby: Be sure to get out and vote in this key election in our country! I did!!! #ivotedtoday #ElectionNight #Elections2016 @77WABC
BaseballBeerBBQ|HappyHourNet|0.7712|0.0|0.691|0.309|RT @HappyHourNet: It's the Nikki X Happy Hour #ElectionDay Special! Tonight at 7:30 ET https://t.co/DyeN4Q0EFY @DrJimmyStar @JETAR9 @LadyLa
BaseballBeerBBQ|blogtalkradio|0.7712|0.0|0.691|0.309|RT @HappyHourNet: It's the Nikki X Happy Hour #ElectionDay Special! Tonight at 7:30 ET https://t.co/DyeN4Q0EFY @DrJimmyStar @JETAR9 @LadyLa
ikkelinear|NewsBud_|-0.5267|0.185|0.815|0.0|RT @NewsBud_: Did Russia Hack the Election? A Short History of CIA Election Sabotage https://t.co/PK6aTk1V6N (Video) https://t.co/TS0KPC5GA
ikkelinear|newsbud|-0.5267|0.185|0.815|0.0|RT @NewsBud_: Did Russia Hack the Election? A Short History of CIA Election Sabotage https://t.co/PK6aTk1V6N (Video) https://t.co/TS0KPC5GA
kf4bef|SebGorka|0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
kf4bef||0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
thejoepeach|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
thejoepeach|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Vibrantankles|ICMezzo|-0.4215|0.358|0.473|0.169|"@ICMezzo same. Goddamn, this election is like no other, ever..."
SkinbyKimH|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
kodykpelham11|NoleGameday|0.6114|0.0|0.6|0.4|"RT @NoleGameday: Happy election night, #Noles!  https://t.co/gqzEAWdsDW"
kodykpelham11|twitter|0.6114|0.0|0.6|0.4|"RT @NoleGameday: Happy election night, #Noles!  https://t.co/gqzEAWdsDW"
MxHarperion|blogdiva|0.0|0.0|1.0|0.0|RT @blogdiva: THIS REMINDS ME... are we getting taco trucks on every corner the day after the election or the day after inauguration? #Ele
wawzxz|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
wawzxz|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
ChickWithKicksz|cruzzz_1|0.0|0.0|1.0|0.0|RT @cruzzz_1: I ain't even tryna watch the election today
pauldrawdy|TheBabylonBee|0.0258|0.138|0.718|0.144|"RT @TheBabylonBee: The True Election Was In Eternity Past, Annoying Calvinist Keeps Reminding Everyone https://t.co/IGCNuFrJxL https://t."
pauldrawdy|babylonbee|0.0258|0.138|0.718|0.144|"RT @TheBabylonBee: The True Election Was In Eternity Past, Annoying Calvinist Keeps Reminding Everyone https://t.co/IGCNuFrJxL https://t."
rosie_apperleyy|RLong_Bailey|-0.5|0.177|0.823|0.0|RT @RLong_Bailey: 3 little bits of bad news the Tories slipped out on US Election Day https://t.co/mRHjfhTCkt
rosie_apperleyy|mirror|-0.5|0.177|0.823|0.0|RT @RLong_Bailey: 3 little bits of bad news the Tories slipped out on US Election Day https://t.co/mRHjfhTCkt
starmonkey4304|michaelianblack|-0.0516|0.132|0.746|0.123|RT @michaelianblack: Quick reminder that Paul Ryan and nearly the entire Republican leadership disgraced themselves at every opportunity th
sinfulweeknd|khairounaaaaa|0.3597|0.0|0.889|0.111|"RT @khairounaaaaa: this whole election has shown me how capitalism is a fucking joke, so who's gonna teach me about communism? https://t.co"
sinfulweeknd|t|0.3597|0.0|0.889|0.111|"RT @khairounaaaaa: this whole election has shown me how capitalism is a fucking joke, so who's gonna teach me about communism? https://t.co"
mattleising|jmelikidse|0.0|0.0|1.0|0.0|"RT @jmelikidse: Summing up this election year:Red, White and Blew https://t.co/dPuNqr1Xha"
mattleising|twitter|0.0|0.0|1.0|0.0|"RT @jmelikidse: Summing up this election year:Red, White and Blew https://t.co/dPuNqr1Xha"
damngabbiee|ShaanMKhan|0.3182|0.0|0.905|0.095|RT @ShaanMKhan: Our election system is flawed. Water is wet. And you're a genius for realizing it. We get it. Now go vote please.
gkgguy|AliEWentworth|-0.4753|0.279|0.721|0.0|RT @AliEWentworth: Election watching stress eating chocolate cake!  https://t.co/URJ1tL1pzl
gkgguy|twitter|-0.4753|0.279|0.721|0.0|RT @AliEWentworth: Election watching stress eating chocolate cake!  https://t.co/URJ1tL1pzl
ClaudiuIonutes1|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
iamBoozforeal|rudeboyy|0.0772|0.0|0.902|0.098|Video: Common Freestyles About Hillary Clinton &amp; Voting On Election Day  https://t.co/GKLwSuEZI8 https://t.co/3vdRtLdzD4
ValisWatson|HispanicsTrump|0.4374|0.0|0.874|0.126|RT @HispanicsTrump: This election is coming down to the wire. Please if you haven't already get out and vote Trump!! #ElectionDay
ProudfitAsian|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
8skopar|untappd!|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/fyt1hzBlOl #voteforbeer
8skopar|untappd|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/fyt1hzBlOl #voteforbeer
heavehoorg|heave-ho|0.0|0.0|1.0|0.0|"In Philadelphia, rumors give way to an ordinaryelection https://t.co/DtjMlNBlXK"
trustfaIIs|falIawaytyIer|0.4215|0.0|0.823|0.177|RT @falIawaytyIer: attention america this is your official presidential election ballot. vote wisely. #topdebate
SamSteel10|TheLastRefuge2|0.0|0.0|1.0|0.0|RT @TheLastRefuge2: Thread #1  7:00pm Election Results and Discussion https://t.co/dvp9W1yfpJ https://t.co/1kuDOKqQA4
SamSteel10|theconservativetreehouse|0.0|0.0|1.0|0.0|RT @TheLastRefuge2: Thread #1  7:00pm Election Results and Discussion https://t.co/dvp9W1yfpJ https://t.co/1kuDOKqQA4
jjconceptsinc|badwolf303|-0.4215|0.177|0.823|0.0|"RT @badwolf303: Election Day: Voters encounter machine breakdowns, describe intimidation at the polls  https://t.co/B8UY4Or0bx"
jjconceptsinc|washingtonpost|-0.4215|0.177|0.823|0.0|"RT @badwolf303: Election Day: Voters encounter machine breakdowns, describe intimidation at the polls  https://t.co/B8UY4Or0bx"
Lacy_Casper|Klcampbell_7|0.296|0.1|0.708|0.192|"RT @Klcampbell_7: Instead of worrying about the election, just remember that we serve a God that's greater than any past/future president."
_mandytweets|twitter|0.0|0.0|1.0|0.0|I'm literally too afraid to go to sleep because of this election and I'm not even American..#ElectionNight https://t.co/mnFCzKNtjb
Samantha_Ruko|SarahCAndersen|-0.1531|0.086|0.914|0.0|RT @SarahCAndersen: Need to finish tomorrow's comic but the election is messing with my nerves just a LITTLE https://t.co/XjkCcpqXsV
Samantha_Ruko|twitter|-0.1531|0.086|0.914|0.0|RT @SarahCAndersen: Need to finish tomorrow's comic but the election is messing with my nerves just a LITTLE https://t.co/XjkCcpqXsV
rebekahcoffee|darrensands|-0.4215|0.142|0.787|0.071|RT @darrensands: One of the important stories of this election is black organizers who worked to consolidate young black political power po
Sling|biggs_manno|0.5106|0.0|0.858|0.142|@biggs_manno Come check out Sling - We still have all of the channels and you can signup for tonight's free preview https://t.co/wv7dN9zLsu
Sling|blog|0.5106|0.0|0.858|0.142|@biggs_manno Come check out Sling - We still have all of the channels and you can signup for tonight's free preview https://t.co/wv7dN9zLsu
SatansNipss|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
NameLack467|eliselabottcnn|0.0|0.0|1.0|0.0|RT @eliselabottcnn: Election Day 2016: History arrives from @StCollinson @CNNPolitics https://t.co/rtQLGd5XgT
NameLack467|cnn|0.0|0.0|1.0|0.0|RT @eliselabottcnn: Election Day 2016: History arrives from @StCollinson @CNNPolitics https://t.co/rtQLGd5XgT
DanSmailes|realDenaldTrump|-0.0772|0.16|0.727|0.113|RT @realDenaldTrump: I'm proud to say that no living Republican President or Nominee voted for me this election. Also no living sane person
acstar9|_The6thHokage|0.0|0.0|1.0|0.0|RT @_The6thHokage: America After Today's Election https://t.co/SAO8PbE94B
acstar9|twitter|0.0|0.0|1.0|0.0|RT @_The6thHokage: America After Today's Election https://t.co/SAO8PbE94B
Ricolasjersey|thirdeyedshite|0.0|0.0|1.0|0.0|RT @thirdeyedshite: We record right after the election is decided so you know it's about to be fuego take city 
francistill|latimes|0.0|0.0|1.0|0.0|"RT @latimes: Election results are beginning to come in for Indiana, Kentucky and New Hampshire. Here's where it stands so far: https://t.co"
francistill|t|0.0|0.0|1.0|0.0|"RT @latimes: Election results are beginning to come in for Indiana, Kentucky and New Hampshire. Here's where it stands so far: https://t.co"
NTRL_WMN|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
izzyhaen14|AlecPaplham|0.0|0.0|1.0|0.0|RT @AlecPaplham: Realist words I think I have seen all election https://t.co/YMh8fdmfXE
izzyhaen14|twitter|0.0|0.0|1.0|0.0|RT @AlecPaplham: Realist words I think I have seen all election https://t.co/YMh8fdmfXE
Sammmyyy_25|CNN|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
Sammmyyy_25|twitter|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
OwaseyeI|cnn|0.0|0.0|1.0|0.0|"New: Control of Senate, House up for grabs https://t.co/51Yo1M4as3 #follow for more"
GabrielJ_W|See_Em_Play|-0.7579|0.306|0.694|0.0|RT @See_Em_Play: people to blame if the democrats lose the election: democratsnot to blame: bernie sanders jill stein young people
questiontheLaw|scotthortonshow|0.0|0.0|1.0|0.0|RT @scotthortonshow: Election Night Live Stream https://t.co/OdbsCg7xgw #tlot @LibertarianInst
questiontheLaw|libertarianinstitute|0.0|0.0|1.0|0.0|RT @scotthortonshow: Election Night Live Stream https://t.co/OdbsCg7xgw #tlot @LibertarianInst
cai_bou|_ForeverrYOUNG|0.7506|0.0|0.67|0.33|RT @_ForeverrYOUNG: Everybody in they sophisticated bag for Election Day lol I'm not wit it
kanimozhi|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
ReynoldHawthor2|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
silverfemale1|YerberiaCultura|0.862|0.0|0.455|0.545|"RT @YerberiaCultura: Election viewing party, tomorrow! Free BBQ / more :) https://t.co/44moFZlwuz"
silverfemale1|twitter|0.862|0.0|0.455|0.545|"RT @YerberiaCultura: Election viewing party, tomorrow! Free BBQ / more :) https://t.co/44moFZlwuz"
LaneThomaHewitt|TPM|-0.6486|0.338|0.531|0.13|"RT @TPM: LA Times: 1 dead, 3 injured in active shooting in Azusa, California https://t.co/ngSembdKgz https://t.co/otlaiyvDeV"
LaneThomaHewitt|talkingpointsmemo|-0.6486|0.338|0.531|0.13|"RT @TPM: LA Times: 1 dead, 3 injured in active shooting in Azusa, California https://t.co/ngSembdKgz https://t.co/otlaiyvDeV"
teddybear10449|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
ellieisntonline|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
ellieisntonline|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
raychlp|igorvolsky|0.128|0.154|0.677|0.169|RT @igorvolsky: Wild that we're here on Election Eve unsure if one of the candidates will accept defeat and concede for the good of our dem
ThinkBigGoLocal|instagram|0.0|0.0|1.0|0.0|Voted  Glass of Wine  Waiting on election results  as a #woman #businessowner or #entre https://t.co/yfDnqoeiOZ https://t.co/amlacEfH6B
greenspank|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
greenspank|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
XRoads003|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
XRoads003|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
luletobe|Bohoover|-0.4019|0.144|0.856|0.0|"RT @Bohoover: Utah: Voting Machine Problems Could Force 52,000 to Use Paper Ballots - Breitbart https://t.co/udDJIgjh0l via @BreitbartNews"
luletobe|breitbart|-0.4019|0.144|0.856|0.0|"RT @Bohoover: Utah: Voting Machine Problems Could Force 52,000 to Use Paper Ballots - Breitbart https://t.co/udDJIgjh0l via @BreitbartNews"
solavoxdeus|WDFx2EU8|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
solavoxdeus|t|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
Mambear04|BYP_100|0.0|0.0|1.0|0.0|RT @BYP_100: Don't stand for the pettiness at the polls! Call the election protection hotline! https://t.co/AG5xcRUDgB
Mambear04|twitter|0.0|0.0|1.0|0.0|RT @BYP_100: Don't stand for the pettiness at the polls! Call the election protection hotline! https://t.co/AG5xcRUDgB
australian|antfarmer|0.4927|0.0|0.849|0.151|RT @antfarmer: Paul Kelly is very good here on Trump as a vandal and the decline of America ($) https://t.co/ydGRKhuvHc
australian|theaustralian|0.4927|0.0|0.849|0.151|RT @antfarmer: Paul Kelly is very good here on Trump as a vandal and the decline of America ($) https://t.co/ydGRKhuvHc
Hickory_dickery|The_Servant10|-0.3612|0.091|0.909|0.0|RT @The_Servant10: they say the election rigged if trump loses.. same thing my people say when we get pulled over or when we gotta dig anot
moderndanceman|TeamTrump|-0.0772|0.105|0.802|0.093|"RT @TeamTrump: If there's one thing you must share before Election Day, it's this. @realDonaldTrump's closing argument to the American vote"
WesternXTheShow|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
WesternXTheShow|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
marnierussell04|MetalOllie|-0.7845|0.283|0.717|0.0|"RT @MetalOllie: No. This is what is commonly known as an ""election"". One of those things you keep losing, you haunted, frog-faced pissbag."
BeverleeHughes3|benchmarkpol|0.6239|0.0|0.83|0.17|"RT @benchmarkpol: Final prediction: Clinton 87% likely to win, 322 EV to 216. Follow our election coverage tomorrow on twitter! https://t.c"
BeverleeHughes3||0.6239|0.0|0.83|0.17|"RT @benchmarkpol: Final prediction: Clinton 87% likely to win, 322 EV to 216. Follow our election coverage tomorrow on twitter! https://t.c"
dee_mainey|NateSilver538|0.5093|0.0|0.852|0.148|"RT @NateSilver538: Our final forecast of the year just published! Clinton is a 71% favorite in polls-only, 72% in polls-plus. https://t.co/"
dee_mainey|t|0.5093|0.0|0.852|0.148|"RT @NateSilver538: Our final forecast of the year just published! Clinton is a 71% favorite in polls-only, 72% in polls-plus. https://t.co/"
TamaraTattles|CNN|0.0|0.0|1.0|0.0|"@CNN  based in ATLANTA, is suddenly figuring out that we are a very dark shade of pink on this election. I don't think they expected it."
leannelovsin|voguemagazine|0.0|0.0|1.0|0.0|"RT @voguemagazine: ""She doesnt realize it yet, but Election Day is a moment in history for both of us."" https://t.co/aP0pq0q274"
leannelovsin|vogue|0.0|0.0|1.0|0.0|"RT @voguemagazine: ""She doesnt realize it yet, but Election Day is a moment in history for both of us."" https://t.co/aP0pq0q274"
KeswickPinhead|SenFallon2016|0.2481|0.089|0.786|0.125|"RT @SenFallon2016: This election is rigged! I intended to vote for #Trump today, when Jesus smacked me upside the head &amp; made my hand vote"
WeirdWestRadio|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
WeirdWestRadio|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
cmhubbard3446|IngramSmith|0.0|0.0|1.0|0.0|"@IngramSmith @Nolecast ... turns off election coverage and immediately goes to Soundcloud, because priorities."
cskrib94|chrisbharrison|0.0|0.0|1.0|0.0|RT @chrisbharrison: Tonight..in the most dramatic election ever..2 candidates..only one will make it to the White House (read in Harrison v
Chrisrlamar|DTorday|-0.4497|0.235|0.624|0.141|"@DTorday @JamesOKeefeIII @daveweigel but you're cheating the election for Hillary, so how is that fair?"
RainManDigital|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
RainManDigital|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
ScreenplaySnob|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
ScreenplaySnob|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
RM001_Director|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
RM001_Director|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
charprat44|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
charprat44|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
Hernandez_Hates|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
Hernandez_Hates|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
kaylabeight|dana_tonkinson|-0.3818|0.115|0.885|0.0|RT @dana_tonkinson: I don't understand why people are getting upset that people who can't vote are actually getting involved in the electio
FromBactaTank|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
FromBactaTank|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
JakeLapin_syr|NewhouseSports|0.1531|0.0|0.904|0.096|Solid crowd tonight as National Anthem underway on election night here at the Dome @NewhouseSports https://t.co/V1aEpxYm5F
JakeLapin_syr|twitter|0.1531|0.0|0.904|0.096|Solid crowd tonight as National Anthem underway on election night here at the Dome @NewhouseSports https://t.co/V1aEpxYm5F
boezuvsofs|NBCDFW|0.5826|0.0|0.799|0.201|@NBCDFW Election day mammaries ! Thanks for keeping us abreast of the news....what an arresting sight !!
ChiefCRX340|BlastingNews|0.0|0.0|1.0|0.0|RT @BlastingNews: #election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR http
ChiefCRX340|us|0.0|0.0|1.0|0.0|RT @BlastingNews: #election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR http
tiffanysuckkaa|KathleenLights1|0.4199|0.141|0.573|0.286|RT @KathleenLights1: Hope everyone voted today! This election has traumatized me.... I pray for America.
wmarsburg|SusanCalman|0.3612|0.0|0.848|0.152|RT @SusanCalman: Now for the election. I'm staying up all night.  I have provisions. I'm ready.
ContempraINN|HuffPostPol|0.0|0.0|1.0|0.0|These photos of dogs voting are getting us through Election Day https://t.co/oUrkbuPdtE #Endeavor via @HuffPostPol #ElectionDay #Dogs
ContempraINN|huffingtonpost|0.0|0.0|1.0|0.0|These photos of dogs voting are getting us through Election Day https://t.co/oUrkbuPdtE #Endeavor via @HuffPostPol #ElectionDay #Dogs
Huntgolfride|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
terunugah||0.0|0.0|1.0|0.0|come watch the election @ my house!
BrooklynnRamos|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
BrooklynnRamos|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
CEntertainment3|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
CEntertainment3|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
CrossroadsSPN|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
CrossroadsSPN|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
DConCW|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
DConCW|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
CritiqueRevolve|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
CritiqueRevolve|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
greeneyes3855|twitter|0.4019|0.0|0.895|0.105|"Though this Election has brought out my PTSD I know I do not stand alone,I WILL NOT BE TAKING RX MEDS to help me th https://t.co/jyK0pgf9Fu"
CazadorProd|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
CazadorProd|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
CeeStormborn|barstoolsports|0.5719|0.0|0.856|0.144|"RT @barstoolsports: Before you move to Canada after this election, learn some more about our neighbors to the north. They're happy to have"
ASixGunForLobo|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
ASixGunForLobo|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
dericdunk|mike_pence|0.3818|0.0|0.894|0.106|"RT @mike_pence: The outcome of this historic election rests in your hands. If you stand for a stronger America, cast your vote for #TrumpPe"
poooyak|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
poooyak|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
gc_wilson|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
novembereve|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
PatriotIBRWB|RealDJTrumpTeam|0.2124|0.0|0.934|0.066|"RT @RealDJTrumpTeam: Don't let up, get out to vote - this election is FAR FROM OVER! We are doing well but there is much time left. GO #FLO"
Okavangomick|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
Okavangomick|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
Mrgee_bande|Telegraph|0.0|0.0|1.0|0.0|RT @Telegraph: Florida polls start closing in less than 10 minutes. It's a crucial state to watch on #ElectionNight https://t.co/CJCBsKKKNE
Mrgee_bande|telegraph|0.0|0.0|1.0|0.0|RT @Telegraph: Florida polls start closing in less than 10 minutes. It's a crucial state to watch on #ElectionNight https://t.co/CJCBsKKKNE
coldplayitcool|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
coldplayitcool|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
jwbrower|twitter|0.6588|0.0|0.672|0.328|Election pizza is so '90s. The #ElectionChili is great! https://t.co/Fsy4nLs9mX
cmdr_hellstorm|twitter|0.1779|0.173|0.578|0.249|Just in case Hilary wins the election and a war really breaks out with Russia ;) https://t.co/83ktE2OWeM
__gacissej|tbhjuststop|0.6249|0.0|0.661|0.339|RT @tbhjuststop: A great way to start Election Day https://t.co/2G8kT6ZyuE
__gacissej|twitter|0.6249|0.0|0.661|0.339|RT @tbhjuststop: A great way to start Election Day https://t.co/2G8kT6ZyuE
miracles3337|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
miracles3337||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
KaylaNoe1|WORLDSTAR|0.5859|0.0|0.678|0.322|RT @WORLDSTAR: Who will win the 2016 presidential election? 
AngelaTGregory|WAVY_News|0.0|0.0|1.0|0.0|Polls are about to close in Virginia. Watch @WAVY_News for complete election results. #Election2016
steve62269|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
INFOS_EN|belfasttelegraph|0.25|0.0|0.824|0.176|US election results: Donald Trump and Hillary Clinton await their verdict of voters - Belfast Telegraph https://t.co/ypMwah7jqC
theNeutral00|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
theNeutral00|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
arembooks|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
arembooks|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
Bamboy360|timkmak|0.3182|0.0|0.897|0.103|RT @timkmak: 4Chan on Election Day Maybe next time try getting an actual competent politician as a nominee instead of a meme. https://t.c
Bamboy360||0.3182|0.0|0.897|0.103|RT @timkmak: 4Chan on Election Day Maybe next time try getting an actual competent politician as a nominee instead of a meme. https://t.c
lissxette|DarkerThanAkon|0.0|0.0|1.0|0.0|RT @DarkerThanAkon: IT'S ELECTION DAY I KNOW YA'LL WILL MAKE THE RIGHT DECISION https://t.co/yF73IzfIk4
lissxette|twitter|0.0|0.0|1.0|0.0|RT @DarkerThanAkon: IT'S ELECTION DAY I KNOW YA'LL WILL MAKE THE RIGHT DECISION https://t.co/yF73IzfIk4
MrFijiWiji|VentureDZN|0.0|0.0|1.0|0.0|RT @VentureDZN: Remember to vote for @MrFijiWiji this election #PutABigBoyIncharge
aeoost|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
aeoost|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
BrooksLandgraf|WillHurd|0.4574|0.0|0.834|0.166|RT @WillHurd: WATCH: Special Election Day Message from Will Hurd! #TX23 #KeepTexasRedFor polling information visit: https://t.co/BgwhQTaM
BrooksLandgraf|t|0.4574|0.0|0.834|0.166|RT @WillHurd: WATCH: Special Election Day Message from Will Hurd! #TX23 #KeepTexasRedFor polling information visit: https://t.co/BgwhQTaM
increase32|TravisRuger|-0.2263|0.203|0.642|0.155|RT @TravisRuger: A vote for Hillary is supporting election fraud.    #PodestaEmails33 #ElectionFinalThoughts #DNCLeaks2 #NeverHillary https
lucidglitch|meakoopa|0.0|0.0|1.0|0.0|"RT @meakoopa: this election I learned a lot about liberalism and the word ""we."" https://t.co/M6wUoce9G5"
lucidglitch|twitter|0.0|0.0|1.0|0.0|"RT @meakoopa: this election I learned a lot about liberalism and the word ""we."" https://t.co/M6wUoce9G5"
villarreal1375|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
kssturgeon|KOINCurt|0.0|0.0|1.0|0.0|RT @KOINCurt: Election night for journalists. @JournalistsLike https://t.co/p6vm8ctjTp
kssturgeon|twitter|0.0|0.0|1.0|0.0|RT @KOINCurt: Election night for journalists. @JournalistsLike https://t.co/p6vm8ctjTp
BBC|BBCWorld|0.1695|0.0|0.894|0.106|RT @BBCWorld: Follow @BBCUSElection for #ElectionNight results &amp; our ongoing coverage &amp; analysishttps://t.co/HkEjD3a3YG*don't forget co
BrockPolly|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
XiamenSec|yahoo|0.0|0.0|1.0|0.0|Stock futures tick up ahead of U.S. election results: https://t.co/I6hrjBQbxn
PA_to_SoCal|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
itznick2|MattZupon|0.0|0.0|1.0|0.0|RT @MattZupon: See my 2016 presidential prediction map |  https://t.co/T9HLo4qHOA
itznick2|foxnews|0.0|0.0|1.0|0.0|RT @MattZupon: See my 2016 presidential prediction map |  https://t.co/T9HLo4qHOA
FearDept|CharlotteHall26|-0.4404|0.153|0.847|0.0|RT @CharlotteHall26: I'm scared for this election result come on America make the right choice  #ElectionNight https://t.co/YMWR6Zfebt
FearDept|twitter|-0.4404|0.153|0.847|0.0|RT @CharlotteHall26: I'm scared for this election result come on America make the right choice  #ElectionNight https://t.co/YMWR6Zfebt
Sovual|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
_tieeee|twitter|0.0|0.0|1.0|0.0|"With this election, YALL DONT HAVE MUCH TIME https://t.co/MXA9qkWxxh"
Waja1130|kmbiamnozie|0.0|0.0|1.0|0.0|"RT @kmbiamnozie: An estimated 150,000 Haitian-American voters live in Florida, the state where 537 votes decided the 2000 election, Trump"
lappinm|tancredipalmeri|0.7901|0.0|0.696|0.304|@tancredipalmeri This is the superb Jeremy Vine! Election maestro extraordinaire who helps us make sense of it all.
LucyTheKhaleesi|twitter|0.0|0.0|1.0|0.0|This election https://t.co/GSQxhMgUzq
acottos|twitter|0.6884|0.12|0.559|0.321|Students participated in a mock election today! Great civics lesson! Thank you students for your participation! https://t.co/R3AmWkZtRy
Kiajanae23|__Shaquille__|-0.5927|0.181|0.75|0.069|RT @__Shaquille__: I'm ready for this election to be over...it's not doing anything but revealing how stupid n uneducated some people are..
CellarDoorSkep|PaleoRadioShow|0.0|0.0|1.0|0.0|"RT @PaleoRadioShow: Our #FinalElectionThoughts on #Election2016, @Wikileaks &amp; future of MSM, and PaleoRadio's role in #atheist punditry! ht"
ihearthestia|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
jamhow2|HuffingtonPost|0.0|0.0|1.0|0.0|RT @HuffingtonPost: 30 oddly insightful quotes from kids about the election https://t.co/0WwtoflHHU https://t.co/2ghyhcKAOh
jamhow2|m|0.0|0.0|1.0|0.0|RT @HuffingtonPost: 30 oddly insightful quotes from kids about the election https://t.co/0WwtoflHHU https://t.co/2ghyhcKAOh
arctic_glitch|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
Lermont|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
kadar_k|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
kadar_k|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
a7xrocker1981|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you VOTED TO DRAIN THE SWAMP! #MAGA #ElectionDay #Election https://t.co/TkUPGBNYkg
a7xrocker1981|twitter|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you VOTED TO DRAIN THE SWAMP! #MAGA #ElectionDay #Election https://t.co/TkUPGBNYkg
tamaraleighllc|RickRWells|0.0772|0.133|0.718|0.149|RT @RickRWells: Has Valerie Jarrett Convinced Obama To Fire Comey After The Election? https://t.co/VmVUcK1zo5 https://t.co/MwlM7UkrKY
tamaraleighllc|stopthetakeover|0.0772|0.133|0.718|0.149|RT @RickRWells: Has Valerie Jarrett Convinced Obama To Fire Comey After The Election? https://t.co/VmVUcK1zo5 https://t.co/MwlM7UkrKY
HabDestini|HabPria|-0.296|0.121|0.879|0.0|Why is @HabPria telling who should have an opinion on a #Election? You're no Barack Obama babes... Xo
seminary_bros|BYUSportsNation|-0.4588|0.167|0.833|0.0|"RT @BYUSportsNation: #BYUSN Election Day Poll - Proposition 3Should the word ""ELITE"" be banned from @Spencer_Linton's vocabulary?"
NajetteDhabi|channeltennews|0.0|0.0|1.0|0.0|RT @channeltennews: #BREAKING: Reports 4 people wounded after shooting near a polling station in Azusa California. #TenNews https://t.co/O0
NajetteDhabi|t|0.0|0.0|1.0|0.0|RT @channeltennews: #BREAKING: Reports 4 people wounded after shooting near a polling station in Azusa California. #TenNews https://t.co/O0
TrentJarrod|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
hapinachu|IZOD|0.296|0.0|0.804|0.196|RT @IZOD: Election Day. Share your voice with #MyVote2016 https://t.co/IDvaKYOxxy
hapinachu|twitter|0.296|0.0|0.804|0.196|RT @IZOD: Election Day. Share your voice with #MyVote2016 https://t.co/IDvaKYOxxy
SnoVitKatt|livsiegfried|0.0|0.0|1.0|0.0|RT @livsiegfried: Looking forward to staying up and watching the election with @TheYoungTurks #tytlive #ElectionDay #ElectionNight https://
SnoVitKatt||0.0|0.0|1.0|0.0|RT @livsiegfried: Looking forward to staying up and watching the election with @TheYoungTurks #tytlive #ElectionDay #ElectionNight https://
peggy_fruge|SebGorka|0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
peggy_fruge||0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
HildaG75|Chrisdr504|0.0|0.0|1.0|0.0|RT @Chrisdr504: May the election night drinking commence! https://t.co/6lhiSTXDK7
HildaG75|twitter|0.0|0.0|1.0|0.0|RT @Chrisdr504: May the election night drinking commence! https://t.co/6lhiSTXDK7
jane9668|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
Michaelcraddo16|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Beto10cafetero|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Beto10cafetero|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
FayForever_|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
FayForever_|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
peachgrI|pupbasket|0.5719|0.0|0.821|0.179|RT @pupbasket: If Trump   Wins The Election I Am Moving   Out Of The Country  Goodbye   America   Hello   EXO Planet 
WillRowland7|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
kimmurphy|latimes|0.0|0.0|1.0|0.0|Exit polls: white college-educated voters trending more Democrat than 2012. Non-college educated whites? Trump town. https://t.co/u0nbNhr8ee
ustadhizmeteri|DahiBilal|0.0|0.0|1.0|0.0|@DahiBilal @TayyipAga Sayin @realDonaldTrump  ve @HillaryClinton This is election result from Usa so far according to @ahbrtv
ericwormann|ConAirFan|0.0772|0.108|0.772|0.12|"RT @ConAirFan: Media tries to discourage voting by dropping ""John Lithgow was originally cast as Frasier on Cheers"" story on election eve."
rcbbstcrk|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
berlinbarbarism|thebafflermag|0.0|0.0|1.0|0.0|RT @thebafflermag: Journalists have been far more attentive to their racial biases than their class biases this election cycle. https://t.c
berlinbarbarism||0.0|0.0|1.0|0.0|RT @thebafflermag: Journalists have been far more attentive to their racial biases than their class biases this election cycle. https://t.c
IsaHerrera_8|latimes|0.0|0.0|1.0|0.0|"RT @latimes: Election results are beginning to come in for Indiana, Kentucky and New Hampshire. Here's where it stands so far: https://t.co"
IsaHerrera_8|t|0.0|0.0|1.0|0.0|"RT @latimes: Election results are beginning to come in for Indiana, Kentucky and New Hampshire. Here's where it stands so far: https://t.co"
diiks_|AmandaPBernard|0.296|0.0|0.732|0.268|RT @AmandaPBernard: This election is a joke #ElectionNight
Suweetpea|FredZeppelin12|0.25|0.0|0.895|0.105|RT @FredZeppelin12: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERS. Advantage #Trump. Evening voters are evening voters because t
YawNinno|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
YawNinno|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
CarloJose1718|ThomasMeikrantz|0.0|0.0|1.0|0.0|That's why meanwhile @ThomasMeikrantz tell me any developments on Salisbury High School girls soccer vs Montoursville and @NBCNews election
tlvrp_russia|therussophile|-0.3818|0.157|0.843|0.0|#Moscow #SaintPetersburg WikiLeaks must publish and be damned: Assange address on US election day https://t.co/OOTNnQ0YoC
MsLake1|dailycal|0.0|0.0|1.0|0.0|Election night drinking game | The Daily Californian https://t.co/EpsUU4YlVQ
XtarTalk|politico|0.3612|0.0|0.762|0.238|How to watch Election Day like a pro https://t.co/gr5T7iRVVU #election2016
jazminxrod|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: Florida, its Election Day! Polls are open from 7am-7pm. Confirm your polling place now and go vote for Hillary! https:"
Magic_C123|Things4WhitePpl|0.0|0.0|1.0|0.0|"""@Things4WhitePpl: Breaking up over an election. https://t.co/du9QC9NaG2"""
Magic_C123|twitter|0.0|0.0|1.0|0.0|"""@Things4WhitePpl: Breaking up over an election. https://t.co/du9QC9NaG2"""
ThatJaysFan20|CJR16255|0.0|0.0|1.0|0.0|"@CJR16255 are you talking about the election or the gold gloves, etc? because I'm ineligible to vote for either"
travis_switala|ayyitsDolan|-0.8381|0.42|0.58|0.0|"RT @ayyitsDolan: I hate politics, I can't wait for this shitty election to be over"
raincoaster|5150committee|-0.7856|0.284|0.716|0.0|"RT @5150committee: It's not clear yet how this election is going to turn out, but what is clear is that it's @Snowden's fault."
Matthanks1|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Matthanks1|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
jensenoliviaa|twitter|0.6696|0.0|0.71|0.29|the best episode of gilmore girls to watch on election day! https://t.co/043P6u5lgg
HiImSerenity|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
HiImSerenity|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
Andrew_Tuft|TBNSport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
Andrew_Tuft|tbnsport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
allie_renee11|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
snipermoney412|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
snipermoney412|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
bushi_jp|youtube|0.0|0.0|1.0|0.0|"""USA: New Yorkers face long queues as they cast their votes in 2016 US election""  YouTube  https://t.co/cpyYnnkmLk"
thedestgroup|realtor|0.6052|0.0|0.78|0.22|Election? What Election?! Check Out These Cute Animals We Found in Listing Photos! https://t.co/EPMnWfskDU https://t.co/eri8sHuXL9
SAILORSOLEMN|CNNPolitics|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
SAILORSOLEMN|twitter|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
XiamenSec|yahoo|0.0|0.0|1.0|0.0|Futures tick up ahead of U.S. election results: https://t.co/ZY3bRZsEuu
patnaikanu|VP|0.0|0.0|1.0|0.0|RT @VP: Today is Election Day in America. Its time to get out and vote. https://t.co/a0MJUF4QIy
patnaikanu|twitter|0.0|0.0|1.0|0.0|RT @VP: Today is Election Day in America. Its time to get out and vote. https://t.co/a0MJUF4QIy
kmsangelica|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
kmsangelica|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
INFOS_EN|bustle|0.4019|0.0|0.838|0.162|"""Pantsuit Nation"" Stories About Voting For Hillary Clinton Offer A Home Stretch Election Boost - Bustle https://t.co/XFy9b3f4WW"
rileeeees|VeronicaRuckh|-0.0653|0.099|0.774|0.128|"RT @VeronicaRuckh: TBH the worst thing about this election is the ""vote shaming."" Everyone's like ""it's so important that you vote,"" but th"
GetSetGoBand|twitch|0.4522|0.0|0.859|0.141|"So, I'm doing a special Election Night show this evening. The pre-show starts at 6:00pm Central (in two minutes.)... https://t.co/Kn6TBNKySj"
EricFreckman|instagram|0.0|0.0|1.0|0.0|Election Day  https://t.co/EDcwdtMf8G
RoxerSoDevious|InappropriateSB|0.0|0.0|1.0|0.0|RT @InappropriateSB: This election in a nutshell https://t.co/TE1m8Scmmi
RoxerSoDevious|twitter|0.0|0.0|1.0|0.0|RT @InappropriateSB: This election in a nutshell https://t.co/TE1m8Scmmi
douglasIsles|youtube|0.4019|0.0|0.803|0.197|Expect #Beyonc to receive to royalty boost as election results announced : https://t.co/G2O2QOpebH
brittan60903516|BaeFeeling|0.0|0.0|1.0|0.0|RT @BaeFeeling: Twitter on Election Day https://t.co/YOLTWcDeqN
brittan60903516|vine|0.0|0.0|1.0|0.0|RT @BaeFeeling: Twitter on Election Day https://t.co/YOLTWcDeqN
BethB1213|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
BethB1213||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
Allypapa_|B96Chicago|0.0|0.0|1.0|0.0|RT @B96Chicago: . @FifthHarmony's @camilacabello97 on #Election2016: 'Immigration is What This Country was Built On' https://t.co/kxfcWoIfd
Allypapa_|t|0.0|0.0|1.0|0.0|RT @B96Chicago: . @FifthHarmony's @camilacabello97 on #Election2016: 'Immigration is What This Country was Built On' https://t.co/kxfcWoIfd
uzzi24|DavidShuster|0.5423|0.0|0.791|0.209|"RT @DavidShuster: Weather channel until 12am:  ""escape the election:  marathon to evoke tranquility, featuring weather scenes set to a rela"
Juan_Migg|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
Juan_Migg|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
kmcfadzen|BrundageKV|0.0|0.0|1.0|0.0|RT @BrundageKV: SAS Elementary students watching US election results in ES Library! #sasedu #USElection2016 https://t.co/OU03Okb4Sa
kmcfadzen|twitter|0.0|0.0|1.0|0.0|RT @BrundageKV: SAS Elementary students watching US election results in ES Library! #sasedu #USElection2016 https://t.co/OU03Okb4Sa
andregreen0|CNN|0.6369|0.0|0.833|0.167|"RT @CNN: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/QurbNzL1BK"
andregreen0|cnn|0.6369|0.0|0.833|0.167|"RT @CNN: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/QurbNzL1BK"
RyanRMiner|twitter|0.0|0.0|1.0|0.0|Which website will you be using for real-time election results. https://t.co/uEWek0ra6W
NotcoolOToole|TheTrumpPuppet|0.0|0.0|1.0|0.0|"RT @TheTrumpPuppet: ""Hello Hillary. How are you doing?"" #Trump #TheTrumpPuppet #Election #ElectionDay https://t.co/iPeB6nFXbl"
NotcoolOToole|vine|0.0|0.0|1.0|0.0|"RT @TheTrumpPuppet: ""Hello Hillary. How are you doing?"" #Trump #TheTrumpPuppet #Election #ElectionDay https://t.co/iPeB6nFXbl"
PencilShank|wired|0.0|0.0|1.0|0.0|Watch WIRED and Ozys Election Night Livestream - https://t.co/FfWqINZ0Qk https://t.co/vXtMOxbwm7
Richard_RSC|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
Richard_RSC|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
HIGHLYBISEXUAL|THOTJAI|0.5719|0.0|0.821|0.179|RT @THOTJAI: if donald trump wins the election I will paypal 100 dollars to everyone that retweets this #ElectionDay
ShaneGasiorows1|HIGH_TIMES_Mag|0.2225|0.0|0.921|0.079|RT @HIGH_TIMES_Mag: We're back on FB Live! Want to know the second weed gets legalized? IGH TIMES is covering the election live! https://t.
ShaneGasiorows1||0.2225|0.0|0.921|0.079|RT @HIGH_TIMES_Mag: We're back on FB Live! Want to know the second weed gets legalized? IGH TIMES is covering the election live! https://t.
Leandra_C_Lee|lntroset|0.8969|0.0|0.67|0.33|RT @lntroset: Today is Election Day so I thought I would share the loving someone lyrics with you guys bc this world needs more love and le
Refinery29|refinery29|0.4588|0.0|0.75|0.25|How your favorite celebs are voting during #ElectionDay: https://t.co/OWRZ0dyO0m https://t.co/OyC6vTclZ9
YesOrMo|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
YesOrMo|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
GladIsLovinNews|business|0.0|0.0|1.0|0.0|RT @business: Both candidates went to the polls this morning in New York https://t.co/MWmkuavh72 #ElectionNight https://t.co/8p58SdCge9
GladIsLovinNews|bloomberg|0.0|0.0|1.0|0.0|RT @business: Both candidates went to the polls this morning in New York https://t.co/MWmkuavh72 #ElectionNight https://t.co/8p58SdCge9
TheMassesAwaken|vefanturmandos|0.6808|0.0|0.741|0.259|"@vefanturmandos @mitchellvii Good to hear. Yes, this election won't be over for another day or two at least."
ideep9|theverge|0.0|0.0|1.0|0.0|verge: 10 provocative political novels to read after the election https://t.co/GW4jdHfTae  https://t.co/l3B4bwr5qC
sean_r_moore|"lerdody,"|0.6696|0.0|0.71|0.29|"Follow @lerdody, @hayleighcolombo, and @IBJnews for the best election coverage tonight! https://t.co/sF1dG2uKIt"
sean_r_moore|twitter|0.6696|0.0|0.71|0.29|"Follow @lerdody, @hayleighcolombo, and @IBJnews for the best election coverage tonight! https://t.co/sF1dG2uKIt"
AuburnFox11|Bencjacobs|0.0|0.0|1.0|0.0|RT @Bencjacobs: Cash bar at trump election night event
MattMaaisas|Jonbuckhouse|0.6239|0.0|0.843|0.157|RT @Jonbuckhouse: The Polls are starting to close all over the US! Who do you think will win the election?  #ElectionNight #electionday #iV
90sBabyTay|BIackPplVids|0.5719|0.0|0.748|0.252|RT @BIackPplVids: Back in 2012 when Obama won the 2012 election  https://t.co/nvEENKBnqj
90sBabyTay|twitter|0.5719|0.0|0.748|0.252|RT @BIackPplVids: Back in 2012 when Obama won the 2012 election  https://t.co/nvEENKBnqj
izzzz22|sports|0.0|0.0|1.0|0.0|LmaoRic Flair voted for Ric Flair for president https://t.co/G1f1zNaXed
jrwsjs|recordonline|0.4404|0.0|0.847|0.153|RT @recordonline: Here's what Trump and Clinton supporters are saying about this historic Election Night https://t.co/lgWpBu129k https://t.
jrwsjs|recordonline|0.4404|0.0|0.847|0.153|RT @recordonline: Here's what Trump and Clinton supporters are saying about this historic Election Night https://t.co/lgWpBu129k https://t.
_michellehinman|Arianaajpg|-0.6124|0.211|0.789|0.0|RT @Arianaajpg: this election has brought out all the racist people that still exist in America...sad
kodykpelham11|astrick005|0.7579|0.082|0.648|0.27|RT @astrick005: Just had someone in verizon argue with me that whoever wins the election immediately goes into office tomorrow I love worki
potential5661|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: Drudge saying, ""Election will come down to evening voters.""  That means, ""Republicans with actual jobs."""
OohNina|janeosanders|0.6369|0.071|0.66|0.269|"RT @janeosanders: Nice story &amp; video re: our incredible supporters  tough day, various choices. #OurRevolution endures. https://t.co/E6Vbi"
OohNina|t|0.6369|0.071|0.66|0.269|"RT @janeosanders: Nice story &amp; video re: our incredible supporters  tough day, various choices. #OurRevolution endures. https://t.co/E6Vbi"
dubhlann123|anne_theriault|0.0|0.0|1.0|0.0|@anne_theriault You can't buy alcohol on election day in Indiana!  *sob*
AlicePolidoro|surfermom77|0.0|0.0|1.0|0.0|"RT @surfermom77: Twitter &amp; FB R begin inundated wt reports of Elec.fraud, voting irregularities &amp; discrimination against Trump Votershttps"
Makaola|inHERribs|0.0|0.0|1.0|0.0|RT @inHERribs: Election Day.  https://t.co/iCYTjRIbn4
Makaola|twitter|0.0|0.0|1.0|0.0|RT @inHERribs: Election Day.  https://t.co/iCYTjRIbn4
BillWestbrook|Franklin_Graham|0.765|0.0|0.714|0.286|RT @Franklin_Graham: This election isnt overits going to be a tight race. Join with family or friends to pray throughout the night that
mommags2579|_IAmChrono_|0.5859|0.0|0.678|0.322|RT @_IAmChrono_: Who should win this election ? #myvote2016   #ElectionDay
JocyTorralba|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
JocyTorralba|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
fifa15sniper123|NBCNews|0.0|0.0|1.0|0.0|"RT @NBCNews: It's just minutes until polls close in Georgia, Indiana, Kentucky, South Carolina, Vermont &amp; Virginia. Follow here: https://t."
fifa15sniper123||0.0|0.0|1.0|0.0|"RT @NBCNews: It's just minutes until polls close in Georgia, Indiana, Kentucky, South Carolina, Vermont &amp; Virginia. Follow here: https://t."
sunday_quilter|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
sunday_quilter||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
Phillygr8|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
TRINITYPRAISE|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
justwaldrop|WalshFreedom|-0.7876|0.338|0.558|0.104|"RT @WalshFreedom: I'm not saying this ELECTION is rigged, but Trump is right: The SYSTEM is rigged. Rigged to help Elites and rigged to s"
garrettrow|shaunna_jayne|0.5719|0.0|0.575|0.425|RT @shaunna_jayne: happy election day  https://t.co/KtwMypK2LL
garrettrow|twitter|0.5719|0.0|0.575|0.425|RT @shaunna_jayne: happy election day  https://t.co/KtwMypK2LL
USA_Votes|usa-votes-2016|0.0|0.0|1.0|0.0|"It's been reported that the LA shooter was ""heavily armed"" https://t.co/7plsFzxyjp #USAVotes2016"
complykated|instagram|0.3612|0.0|0.848|0.152|I remember my parents having election result gatherings. It always seemed like such an adult https://t.co/SwcPUoaP9j
corypheio|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
DarrenjMcLaren|BritishVogue|0.0|0.0|1.0|0.0|RT @BritishVogue: The US Election: What Happens When? https://t.co/sD7EYjbzX3 #ElectionDay https://t.co/ofAJuyfF1k
DarrenjMcLaren|vogue|0.0|0.0|1.0|0.0|RT @BritishVogue: The US Election: What Happens When? https://t.co/sD7EYjbzX3 #ElectionDay https://t.co/ofAJuyfF1k
Marve25|barstoolsports|0.5719|0.0|0.856|0.144|"RT @barstoolsports: Before you move to Canada after this election, learn some more about our neighbors to the north. They're happy to have"
evelynglz_99|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
vampedexo|trapsouIed|0.5719|0.0|0.821|0.179|RT @trapsouIed: If Trump   Wins The Election I Am Moving   Out Of The Country  Goodbye   America   Hello   EXO PLANET
duullcceee_|KeeganAllen|0.6249|0.0|0.843|0.157|"RT @KeeganAllen: Instead of looking at this election as a series finale of the Great American reality show, look at it as your life...start"
explosiveben12|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
explosiveben12|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
WillSmirk4Food|msnbc|-0.4767|0.307|0.693|0.0|"Election night rituals: dinner, porn, crying #maddow https://t.co/5kIlqcnkjv"
Donwood72|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Donald #Trump. Follow @nbcconnecticut for the latest election news.https://t.co/zFdT7UCG1F
coryzsmith|ABC|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
coryzsmith|abcnews|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
ThinkBigGoLocal|facebook|0.0|0.0|1.0|0.0|Voted  Glass of Wine  Waiting on election results  as a #woman #businessowner or #entrepreneur - how concerned... https://t.co/vbMg40OCmk
jamiedelton|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
jamiedelton||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
mite72|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: This election my dad did not spend time raising $ from the billionaire elite. Instead he spent time talking to the Amer
Spicoli83|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
ClarisaS214|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
indystar|AmyBartner|0.0|0.0|1.0|0.0|RT @AmyBartner: We're broadcasting live on https://t.co/gLz3VscwjS with all your live election coverage! https://t.co/NJnVbC4SHZ
indystar|indystar|0.0|0.0|1.0|0.0|RT @AmyBartner: We're broadcasting live on https://t.co/gLz3VscwjS with all your live election coverage! https://t.co/NJnVbC4SHZ
defnii|twitter|-0.4389|0.178|0.724|0.098|This isn't an election! It's a race war against gender started by the MSM and establishment Democrats supported by https://t.co/eVGjagYy9z
sam_rawson96|ZackMUFC|0.7096|0.0|0.685|0.315|"RT @ZackMUFC: Election nights are better than 99% of shite on TV, well worth pulling the all nighter."
andystew22|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
andystew22|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
bjoern_bremer|EconUS|0.0|0.0|1.0|0.0|RT @EconUS: How other countries would vote in the American election https://t.co/noVxb7YGhD https://t.co/Byn4kezRow
bjoern_bremer|economist|0.0|0.0|1.0|0.0|RT @EconUS: How other countries would vote in the American election https://t.co/noVxb7YGhD https://t.co/Byn4kezRow
SirAimnHkim|davidsocomedy|-0.9217|0.41|0.59|0.0|RT @davidsocomedy: P.S.  fuck you dumb fucks hating on anybody tweeting or talking about something other than the election. We all know it'
paulrlanni|GunOwners|-0.6833|0.228|0.772|0.0|RT @GunOwners: Second Amendment rights are literally on the ballot in 5 states. Vote NO on the gun control proposals! #ElectionDay https://
paulrlanni||-0.6833|0.228|0.772|0.0|RT @GunOwners: Second Amendment rights are literally on the ballot in 5 states. Vote NO on the gun control proposals! #ElectionDay https://
kingslayering|dandrego|0.0|0.0|1.0|0.0|"RT @dandrego: can't wait for the election to be over so we can give the polls back to their rightful owners, the strippers"
schwiick|brittanyisbogus|0.8066|0.0|0.644|0.356|"RT @brittanyisbogus: i am feeling very hopeful for this election, hope you all did more than tweet today! https://t.co/TrbkkSEJs5"
schwiick|twitter|0.8066|0.0|0.644|0.356|"RT @brittanyisbogus: i am feeling very hopeful for this election, hope you all did more than tweet today! https://t.co/TrbkkSEJs5"
PattyCamps2|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
KathsBurgess|_KCummings_|0.0|0.0|1.0|0.0|RT @_KCummings_: Election Day 2016 in #JacksonTN. #GoVoteTN https://t.co/LFg7v8D3qn
KathsBurgess|twitter|0.0|0.0|1.0|0.0|RT @_KCummings_: Election Day 2016 in #JacksonTN. #GoVoteTN https://t.co/LFg7v8D3qn
Clintonite33|KellyScaletta|0.4019|0.0|0.856|0.144|"RT @KellyScaletta: ""Active shooter situation"" is NOT something we should see on election day. It's beyond despicable."
envez|cnni|0.0|0.0|1.0|0.0|"RT @cnni: As the 2016 US election campaign ends, follow latest #ElectionNight updates here https://t.co/KMLvpoo10J https://t.co/SRNlKKG6bI"
envez|cnn|0.0|0.0|1.0|0.0|"RT @cnni: As the 2016 US election campaign ends, follow latest #ElectionNight updates here https://t.co/KMLvpoo10J https://t.co/SRNlKKG6bI"
gattacca94|YouTube|0.4215|0.0|0.811|0.189|I liked a @YouTube video https://t.co/E1NQGobAvm USA Election Day 2016 Live - Live Result America Election
gattacca94|youtube|0.4215|0.0|0.811|0.189|I liked a @YouTube video https://t.co/E1NQGobAvm USA Election Day 2016 Live - Live Result America Election
cohnski|vote4wallbanger|0.1027|0.0|0.851|0.149|RT @vote4wallbanger: Me as I await the election results.#ElectionDay https://t.co/gNfD5jtN76
cohnski|twitter|0.1027|0.0|0.851|0.149|RT @vote4wallbanger: Me as I await the election results.#ElectionDay https://t.co/gNfD5jtN76
SamSteel10|TheLastRefuge2|0.0|0.0|1.0|0.0|RT @TheLastRefuge2: Thread #1  7:00pm Election Results and Discussion https://t.co/dvp9W1yfpJ https://t.co/n7sKkZRKm8
SamSteel10|theconservativetreehouse|0.0|0.0|1.0|0.0|RT @TheLastRefuge2: Thread #1  7:00pm Election Results and Discussion https://t.co/dvp9W1yfpJ https://t.co/n7sKkZRKm8
BrianaLathon|people|0.5106|0.0|0.837|0.163|RT @people: All the places you can get free food for voting on #ElectionDay https://t.co/dbJdgAY2pQ via @PeopleFood https://t.co/bqvpOmufZO
BrianaLathon|people|0.5106|0.0|0.837|0.163|RT @people: All the places you can get free food for voting on #ElectionDay https://t.co/dbJdgAY2pQ via @PeopleFood https://t.co/bqvpOmufZO
LittleSugar2529|ABC|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
LittleSugar2529|abcnews|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
IndigoHawthorne|ACTBrigitte|0.0|0.0|1.0|0.0|RT @ACTBrigitte: My personal election message #actforamerica #election2016 #neverhillary https://t.co/dPXGLEUkkh
IndigoHawthorne|youtube|0.0|0.0|1.0|0.0|RT @ACTBrigitte: My personal election message #actforamerica #election2016 #neverhillary https://t.co/dPXGLEUkkh
nscrowba|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
nscrowba|t|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
Newsmanjim|CBSThisMorning|0.0|0.0|1.0|0.0|RT @CBSThisMorning: Oh how this map will change. How Election night begins... #CBSElection  https://t.co/SraM591OGV
Newsmanjim|twitter|0.0|0.0|1.0|0.0|RT @CBSThisMorning: Oh how this map will change. How Election night begins... #CBSElection  https://t.co/SraM591OGV
andrialisa24|chrislhayes|-0.5256|0.159|0.841|0.0|RT @chrislhayes: Trump is already laying the groundwork to contest the legitimacy of the election and it's incredibly dangerous.
jrwsjs|recordonline|0.1027|0.112|0.759|0.129|RT @recordonline: Trump spent a good portion of Election Day sowing doubt about the legitimacy of the election results https://t.co/zdp7B41
jrwsjs|t|0.1027|0.112|0.759|0.129|RT @recordonline: Trump spent a good portion of Election Day sowing doubt about the legitimacy of the election results https://t.co/zdp7B41
amieabenth|swastvedt|0.4574|0.0|0.864|0.136|"RT @swastvedt: You, yes YOU can still register to #Vote2016 in MN! https://t.co/cxQYlNEhSi. More at 11 on @MPRnews w/ @webertom1"
amieabenth|sos|0.4574|0.0|0.864|0.136|"RT @swastvedt: You, yes YOU can still register to #Vote2016 in MN! https://t.co/cxQYlNEhSi. More at 11 on @MPRnews w/ @webertom1"
Leifinator|SarahCAndersen|-0.1531|0.086|0.914|0.0|RT @SarahCAndersen: Need to finish tomorrow's comic but the election is messing with my nerves just a LITTLE https://t.co/XjkCcpqXsV
Leifinator|twitter|-0.1531|0.086|0.914|0.0|RT @SarahCAndersen: Need to finish tomorrow's comic but the election is messing with my nerves just a LITTLE https://t.co/XjkCcpqXsV
woda01|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
woda01|t|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
thatkindofplace|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
Kmpcool123|scumnigger|-0.8047|0.303|0.697|0.0|RT @scumnigger: the election is here but they tryna distract us from the fact childish gambino finna drop his album soon #staywoke
tangopublishing|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
tangopublishing|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
KateSherrill|blogdiva|0.0|0.0|1.0|0.0|RT @blogdiva: THIS REMINDS ME... are we getting taco trucks on every corner the day after the election or the day after inauguration? #Ele
HAYDNRSNAPE|MJosephSheppard|0.7506|0.0|0.701|0.299|RT @MJosephSheppard: Pinellas County Florida Obama won by 5.6 Current two party vote GOP 55% Dem 45%https://t.co/G1z7oNy6Yf
HAYDNRSNAPE|votepinellas|0.7506|0.0|0.701|0.299|RT @MJosephSheppard: Pinellas County Florida Obama won by 5.6 Current two party vote GOP 55% Dem 45%https://t.co/G1z7oNy6Yf
rabuliz|DonaldJTrumpJr|0.3164|0.0|0.906|0.094|RT @DonaldJTrumpJr: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERSGET OUT AND VOTE! Find 5 others. This is our chance to take back Am
len_volkel|shootist2015|0.0|0.0|1.0|0.0|"RT @shootist2015: #Trump smashing #CrookedHillary in early exit poll data from Naples, FL https://t.co/WfaoP82jYN"
len_volkel|naplesnews|0.0|0.0|1.0|0.0|"RT @shootist2015: #Trump smashing #CrookedHillary in early exit poll data from Naples, FL https://t.co/WfaoP82jYN"
Deelishis_Dee|MiamiHerald|0.0|0.0|1.0|0.0|RT @MiamiHerald: Shooting in California leaves two polling places on lock down https://t.co/K46IvO2Mji https://t.co/8pRkf1f2PZ
Deelishis_Dee|miamiherald|0.0|0.0|1.0|0.0|RT @MiamiHerald: Shooting in California leaves two polling places on lock down https://t.co/K46IvO2Mji https://t.co/8pRkf1f2PZ
jvband|AsmSantabarbara|0.1754|0.096|0.783|0.121|"RT @AsmSantabarbara: Proud to cast my ballot in this historic election! If you haven't already, I encourage you to do your part &amp; vote. #El"
Sqwizzey|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
Sqwizzey|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
Wei_Richard|YouTube-Video|0.0|0.0|1.0|0.0|Ich mag das @YouTube-Video: https://t.co/UsWvI2FJ4w Decision 2016: LIVE Election Night Coverage | NBC News
Wei_Richard|youtube|0.0|0.0|1.0|0.0|Ich mag das @YouTube-Video: https://t.co/UsWvI2FJ4w Decision 2016: LIVE Election Night Coverage | NBC News
askhalid|dotlayer8|0.296|0.0|0.833|0.167|"RT @dotlayer8: Surviving 2016: Live election results, memes, and news: https://t.co/2FbMDtlYqa https://t.co/HcLP2wTgLm"
askhalid|dailydot|0.296|0.0|0.833|0.167|"RT @dotlayer8: Surviving 2016: Live election results, memes, and news: https://t.co/2FbMDtlYqa https://t.co/HcLP2wTgLm"
NjdotcomReader|CBCAlerts|0.0|0.18|0.64|0.18|@CBCAlerts Devoting resources to cover another country's election? Probably upsetting a lot of Canadians.
RCRTheRock|TheSweepRU|0.0|0.0|1.0|0.0|Take a break from the election and tune into the @TheSweepRU  in a half hour!
itsyagrlLOLITA|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
itsyagrlLOLITA|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
RenzoNoBenzo_94|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
RenzoNoBenzo_94|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
Klutar|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
Klutar|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
TheShaneHodge|MarianneHaran|0.4199|0.0|0.851|0.149|@MarianneHaran I'll show him what voting 'Other' feels like the next time his is up for election!
PatrickJDuprey|EvanWagstaff|-0.4019|0.144|0.856|0.0|RT @EvanWagstaff: Our #election themed live blog cake. I am that traumatized coder from the second headline https://t.co/3qOFViNC4l
PatrickJDuprey|twitter|-0.4019|0.144|0.856|0.0|RT @EvanWagstaff: Our #election themed live blog cake. I am that traumatized coder from the second headline https://t.co/3qOFViNC4l
CassieMusel|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
atlaswon|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
serina__marie|55mmbae|0.4019|0.0|0.856|0.144|"RT @55mmbae: RT @BreakingNews Independent Party announces new Candidate coming late into the election, Larack Tobama. https://t.co/7ZVTOXiq"
serina__marie|t|0.4019|0.0|0.856|0.144|"RT @55mmbae: RT @BreakingNews Independent Party announces new Candidate coming late into the election, Larack Tobama. https://t.co/7ZVTOXiq"
mmickyon|Reuters|-0.1531|0.118|0.882|0.0|"RT @Reuters: Long lines, raised voices and lawsuits on U.S. #ElectionDay: https://t.co/ulwHwkGMx9 https://t.co/2TIi3XbdC3"
mmickyon|reuters|-0.1531|0.118|0.882|0.0|"RT @Reuters: Long lines, raised voices and lawsuits on U.S. #ElectionDay: https://t.co/ulwHwkGMx9 https://t.co/2TIi3XbdC3"
danshewan|AJemaineClement|0.0|0.0|1.0|0.0|@AJemaineClement he probably understands the election even less than he understood the Brexit vote
mrsmartakis|MattBellassai|-0.0258|0.131|0.742|0.127|"RT @MattBellassai: hey @realDonaldTrump just wanna say that despite everything that's happened this election, you're still awful and i hope"
Avenir078|NPO1|0.0|0.0|1.0|0.0|#electionnight Dutch tv covering the election are too pro #HillaryClinton basically have been talking about her 90% of last hour @NPO1
Andrew__DaSilva|Capitals|0.0|0.0|1.0|0.0|RT @Capitals: When you get to meet a #HoltBeast that's your size. I bet this lil' dude is going to #VoteHoltby. #CapsElectionNight https://
Andrew__DaSilva||0.0|0.0|1.0|0.0|RT @Capitals: When you get to meet a #HoltBeast that's your size. I bet this lil' dude is going to #VoteHoltby. #CapsElectionNight https://
patrickmacsmith|edrummondsmith|0.0|0.0|1.0|0.0|RT @edrummondsmith: Ask a Political Scientist: Election 2016 / Question 5 / White Dudes https://t.co/RAGZFAMAVJ
patrickmacsmith|askapoliticalscientist|0.0|0.0|1.0|0.0|RT @edrummondsmith: Ask a Political Scientist: Election 2016 / Question 5 / White Dudes https://t.co/RAGZFAMAVJ
BeauregardAsher|forctr|0.0|0.0|1.0|0.0|Live updates: Senate election results - https://t.co/QmE1tVMwKs
NotPennn|BrabecNoah|-0.5147|0.322|0.678|0.0|RT @BrabecNoah:  LEAKED RESULTS OF TONIGHT'S ELECTION!  https://t.co/0u8sy9kiZ8
NotPennn|reddit|-0.5147|0.322|0.678|0.0|RT @BrabecNoah:  LEAKED RESULTS OF TONIGHT'S ELECTION!  https://t.co/0u8sy9kiZ8
MynamesJ0y|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
MynamesJ0y|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
freeboy1776|UnifiedPatriots|-0.6486|0.249|0.751|0.0|RT @UnifiedPatriots: from @RealJTP BREAKING: Police Find Texas Election Judge Dead in Home https://t.co/lXzKh0sNhM
freeboy1776|joeforamerica|-0.6486|0.249|0.751|0.0|RT @UnifiedPatriots: from @RealJTP BREAKING: Police Find Texas Election Judge Dead in Home https://t.co/lXzKh0sNhM
Kkowen400Keith|GMA|-0.1027|0.203|0.636|0.161|@GMA at gma your lack of objective reporting and trying to rig election with your hillary favored reports by the minute get ready to suck it
queenbeedrill|ABC|0.0|0.0|1.0|0.0|"RT @ABC: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t.co/Qgyx3"
queenbeedrill|t|0.0|0.0|1.0|0.0|"RT @ABC: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t.co/Qgyx3"
ketch169|seangentille|-0.2714|0.211|0.635|0.154|"RT @seangentille: Thanks to Bill Belichick, you can hate the Patriots again! https://t.co/NlgtjTiwsM https://t.co/vtRDzNeEbf"
ketch169|sportingnews|-0.2714|0.211|0.635|0.154|"RT @seangentille: Thanks to Bill Belichick, you can hate the Patriots again! https://t.co/NlgtjTiwsM https://t.co/vtRDzNeEbf"
BRIMVC|grandelaurminah|0.0|0.0|1.0|0.0|RT @grandelaurminah: We need to make our voices heard for this years election #ImWithHer 
janettwokay|60DaysInFan|0.5719|0.0|0.837|0.163|RT @60DaysInFan: Watching CNN right now and will be watching the whole night to see whom wins The Election. #ElectionNight
PJPsych|cbsnews|0.0|0.0|1.0|0.0|2016 Election Center Live Results - https://t.co/4uUNRYJbJo https://t.co/6VlI53IaJb
david_kennedy11|lolrenaynay|0.4939|0.086|0.703|0.211|"RT @lolrenaynay: Election results come in soon, come here and let me save youFYI I'm drinkingYou can join me, no judgementhttps://t.co/S"
mikeburbachPP|MaraGottfried|0.0|0.0|1.0|0.0|"RT @MaraGottfried: If you're looking for a quick break from election news, here's the story of how Ella Jarman was born on I-94. https://t."
mikeburbachPP||0.0|0.0|1.0|0.0|"RT @MaraGottfried: If you're looking for a quick break from election news, here's the story of how Ella Jarman was born on I-94. https://t."
kristenlongg|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
factiod|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
NASCARNAC|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
WalkerQWalthall|CommonWhiteGrl|0.6249|0.0|0.661|0.339|RT @CommonWhiteGrl: A great way to start Election Day https://t.co/2yM1hzZ36U
WalkerQWalthall|twitter|0.6249|0.0|0.661|0.339|RT @CommonWhiteGrl: A great way to start Election Day https://t.co/2yM1hzZ36U
akepps|tombrokaw.|0.0|0.0|1.0|0.0|Spending my election night with @tombrokaw.  Same as every other presidential election night since I was born.  #NBC #peacock
gissellewbu|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
gissellewbu|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
NCREPUBLICAN|FoxNews|0.0|0.0|1.0|0.0|RT @FoxNews: .@mike_pence &amp; his wife were spotted on a bike ride before the gov. heads to an election center nearby to cast his vote. (VIDE
sydawei|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
GOPbattle2016|mike_pence|0.3818|0.0|0.894|0.106|"RT @mike_pence: The outcome of this historic election rests in your hands. If you stand for a stronger America, cast your vote for #TrumpPe"
alllhypenoheart|BillRatchet|0.765|0.0|0.515|0.485|RT @BillRatchet: i hope whoever wins the election illegalizes anime
M_Jaramillo_333|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
NopeStylinson|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
NopeStylinson|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
louvablesun|armineshaaa|0.0276|0.177|0.641|0.182|RT @armineshaaa: this election is more stressful than that time australia nearly won eurovision https://t.co/jZal4lNpnh
louvablesun|twitter|0.0276|0.177|0.641|0.182|RT @armineshaaa: this election is more stressful than that time australia nearly won eurovision https://t.co/jZal4lNpnh
LeeH3283|ananavarro|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
LeeH3283|twitter|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
OBauby|MsAmyHerron|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
OBauby|theguardian|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
wise_diva|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
wise_diva|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
SadMarchand|dril|0.0|0.0|1.0|0.0|RT @dril: if you ask me this election could end about 100 different ways:1) trump gets 0% of the vote2) trump gets 1% of the vote3) trum
HeyMissHeather|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
HeyMissHeather|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
CANTALINIJON|twitter|-0.3612|0.294|0.706|0.0|Me stressing out about the election: https://t.co/eAztjQjsBF
LoverofAll777|cernovichsdog|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
LoverofAll777|twitter|0.0|0.0|1.0|0.0|RT @cernovichsdog: If I self identify as a human on Election Day - can I vote for Donald J. Trump? #MAGA3X https://t.co/tI8GFaKpxb
jamekiaVsmekia|twitter|0.2411|0.0|0.859|0.141|Election Snack  My decision was with or without nuts  #withnuts #chewies #snacktime https://t.co/dS4ZOiFIjk
msfreakinrosie|jfryer2000|0.0|0.0|1.0|0.0|RT @jfryer2000: Waiting for election results to come in. #ElectionResults #ElectionDay #ElectionNight https://t.co/ZsqleLiTJ3
msfreakinrosie|twitter|0.0|0.0|1.0|0.0|RT @jfryer2000: Waiting for election results to come in. #ElectionResults #ElectionDay #ElectionNight https://t.co/ZsqleLiTJ3
gr00vvyyq|SubMedina|0.0|0.0|1.0|0.0|RT @SubMedina: it's election dayhttps://t.co/IO9qnibSN9
2k_joseph|businessinsider|0.0|0.0|1.0|0.0|RT @businessinsider: LIVE: Results of the 2016 presidential election are rolling in https://t.co/7XwVfYRA6o https://t.co/FOVvXkeF96
2k_joseph|businessinsider|0.0|0.0|1.0|0.0|RT @businessinsider: LIVE: Results of the 2016 presidential election are rolling in https://t.co/7XwVfYRA6o https://t.co/FOVvXkeF96
Halllidisco|tomilo|0.6096|0.0|0.734|0.266|RT @tomilo: This election has given us so many excellent moments... https://t.co/b7SRw2ZIbR
Halllidisco|vine|0.6096|0.0|0.734|0.266|RT @tomilo: This election has given us so many excellent moments... https://t.co/b7SRw2ZIbR
comeandjoinus45|Eileen43Eileen|-0.4019|0.153|0.847|0.0|"RT @Eileen43Eileen: Polling station on lockdown after shooting leaves 4 injured in Azusa, CA  RT America https://t.co/KwZzj2fxBl"
comeandjoinus45|rt|-0.4019|0.153|0.847|0.0|"RT @Eileen43Eileen: Polling station on lockdown after shooting leaves 4 injured in Azusa, CA  RT America https://t.co/KwZzj2fxBl"
SylvieBommel|nytimes|0.5859|0.0|0.787|0.213|"The 1,024 Ways Clinton or Trump Can Win the Election - The New York Times https://t.co/Ake05mmtu6"
Philfandan|BocaRatonRC|0.4404|0.0|0.854|0.146|RT @BocaRatonRC: Who better to torch Hillary to a crisp on election eve than firebrand Tomi Lahren? https://t.co/rnfeyqgAOD https://t.co/4Z
Philfandan|bizpacreview|0.4404|0.0|0.854|0.146|RT @BocaRatonRC: Who better to torch Hillary to a crisp on election eve than firebrand Tomi Lahren? https://t.co/rnfeyqgAOD https://t.co/4Z
MoweryRoger|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Maddman1212|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
ShopTLC007|instagram|0.8698|0.0|0.337|0.663|Happy Election Day!  Almost over! Thank goodness!! https://t.co/kNyASqCzSc
61Rinaldi|hockeydeb21|-0.4466|0.257|0.616|0.128|RT @hockeydeb21: LEAKED CLINTON INTERNAL DOCUMENT: Discourage Trump Supporters with Bogus Polls and Declaring Election Over https://t.co/cJ
61Rinaldi|t|-0.4466|0.257|0.616|0.128|RT @hockeydeb21: LEAKED CLINTON INTERNAL DOCUMENT: Discourage Trump Supporters with Bogus Polls and Declaring Election Over https://t.co/cJ
howelldawson|JoeyGraceffa|0.5461|0.0|0.773|0.227|RT @JoeyGraceffa: RT IF YOU'RE READY FOR THIS ELECTION TO BE OVER!  #ImWithHer
tlvrp_russia|therussophile|0.0|0.0|1.0|0.0|#Moscow #SaintPetersburg Hillary Clinton: A Cabinet Full of Old World Nationalists and Information Operations In C https://t.co/lTgxBfCyzJ
lamaramironova4|cosmopolitan|0.0|0.0|1.0|0.0|Disability-Rights Activist Anastasia Somoza Casts Her Vote for Hillary Clinton https://t.co/r3sZFgLMEi https://t.co/wbjUdkzZyg
Clevohjohn|RussWKYC|-0.5256|0.175|0.825|0.0|@RussWKYC @wkyc @clevelanddotcom very disappointed in the guy I voted for in the primary and the GOV election.
jayoncexomeeka|MASEEZUSWEST|0.0|0.0|1.0|0.0|RT @MASEEZUSWEST: The election effects the whole world soo https://t.co/EcG4osFmCI
jayoncexomeeka|twitter|0.0|0.0|1.0|0.0|RT @MASEEZUSWEST: The election effects the whole world soo https://t.co/EcG4osFmCI
TriXteRPhillips|facebook|0.0|0.0|1.0|0.0|Here is a live stream if you cannot get the Marijuana Election Night 2016 Livestream feed working.... https://t.co/xKMWzwapmk
harpersnotes|projects|0.0|0.0|1.0|0.0|"US election state by state predictions, all one one page. . https://t.co/UHDRJ71nUJ"
BourseetTrading|bloomberg|0.0|0.0|1.0|0.0|#Finance #Trading #Vix keep in mind #ElectionNight https://t.co/G6NN9WUPme https://t.co/lrFuJTfD5e
GoofyNewfie2012|SheldonP|0.0|0.0|1.0|0.0|"@SheldonP Errrmm, USA election night!"
m_abagail|NBCNews|0.296|0.098|0.758|0.144|RT @NBCNews: Can Trump pull an upset in Virginia? The state has been a key to every GOP president's win since 1924: https://t.co/F2MLlKpC7Y
m_abagail|nbcnews|0.296|0.098|0.758|0.144|RT @NBCNews: Can Trump pull an upset in Virginia? The state has been a key to every GOP president's win since 1924: https://t.co/F2MLlKpC7Y
J_Chapz|twitter|0.4215|0.0|0.823|0.177|I've heard stories about election night pizza. I can confirm it's true #electionday  #partylikeajournalist https://t.co/coUyImt4LZ
HillUnfiltered|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
armadillobee|BillRatchet|0.765|0.0|0.515|0.485|RT @BillRatchet: i hope whoever wins the election illegalizes anime
Stella78765322|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
momois|BRANDONWARDELL|0.0|0.0|1.0|0.0|RT @BRANDONWARDELL: election day is peak 4chan https://t.co/AGZkf4PSlN
momois|twitter|0.0|0.0|1.0|0.0|RT @BRANDONWARDELL: election day is peak 4chan https://t.co/AGZkf4PSlN
GunnerLopez|TomBradysEgo|0.7574|0.0|0.629|0.371|RT @TomBradysEgo: Happy Election Day! I think we can all agree on this https://t.co/lxNeiDOp5H
GunnerLopez|twitter|0.7574|0.0|0.629|0.371|RT @TomBradysEgo: Happy Election Day! I think we can all agree on this https://t.co/lxNeiDOp5H
lukey1223|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
aRaymaker|Smaulgld|0.0|0.0|1.0|0.0|RT @Smaulgld: Retweet if you are NOT watching @cnn election coverage tonight
adrianakirk33|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
Hwk765|WalshFreedom|-0.4019|0.351|0.649|0.0|RT @WalshFreedom: Who gives a damn? https://t.co/rJWutS0KlH
Hwk765|thehill|-0.4019|0.351|0.649|0.0|RT @WalshFreedom: Who gives a damn? https://t.co/rJWutS0KlH
CoppedNews|washingtonpost|-0.5859|0.241|0.759|0.0|"#coppednews The Fix: Donald Trump's Election Day insinuations of voter fraud, explained https://t.co/DeLPwh74PL"
LibertVeritJust|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
AbeChristensen|NickTimiraos|0.0|0.0|1.0|0.0|"RT @NickTimiraos: A handy guide to watching election returns: When states to close, and which ones to watch https://t.co/8WPt29yVzb https:/"
AbeChristensen|wsj|0.0|0.0|1.0|0.0|"RT @NickTimiraos: A handy guide to watching election returns: When states to close, and which ones to watch https://t.co/8WPt29yVzb https:/"
tarajoylove|twitter|0.4926|0.0|0.862|0.138|Hope yall got out there &amp; did your part in the most #historic #election ever.  Let them hear us roar! https://t.co/cT0koTTpwi
IvanAlcorchas|biggabossben|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
IvanAlcorchas|twitter|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
LilyDelesse|kbro0ke|0.2023|0.081|0.809|0.11|"RT @kbro0ke: Since no rules are being followed this election season, can we just have four more years of @BarackObama ? He's my fav, anyway."
JooVict18050892|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
ReedG055|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
lunarmuva|benjancewicz|0.0|0.0|1.0|0.0|RT @benjancewicz: Florida voting already surpasses entire 2000 election total https://t.co/DmZLQOG6Sc https://t.co/lzsLjQByup
lunarmuva|cnn|0.0|0.0|1.0|0.0|RT @benjancewicz: Florida voting already surpasses entire 2000 election total https://t.co/DmZLQOG6Sc https://t.co/lzsLjQByup
PlazaRudy|Hardline_Stance|-0.9124|0.493|0.507|0.0|"RT @Hardline_Stance: massive VOTER FRAUD in #FTL #FL; Election workers caught faking 1,000's of stolen absentee ballotshttps://t.co/0ajn3"
Four13Designs|facebook|-0.4019|0.152|0.785|0.063|Escaping the election madness with this prettiness...Hand lettered fabric place cards with a printed topo map of... https://t.co/VRPJ9v0qr5
cuZwersal|miketoews|0.0|0.0|1.0|0.0|@miketoews They'll let you down more than the results of the election...
gandtmilfthree|HotWife937|0.0|0.0|1.0|0.0|RT @HotWife937: HotWifing Election Day    #TittyTuesday #SoMilfy    #MilfieClub #MILFMafia         #RWSW #NGOT           #HotWife h
tjzarro|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
HazaQuiroz|PatrickRothfuss|0.0|0.0|1.0|0.0|RT @PatrickRothfuss: Reminder: In Wisconsin you can register to vote at your polling place on election day.For real. Same-day registratio
frorust|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
Amy12093|IZOD|0.296|0.0|0.833|0.167|RT @IZOD: America votes. Join the Election Day conversation with #MyVote2016 https://t.co/BWuiwAxas6
Amy12093|twitter|0.296|0.0|0.833|0.167|RT @IZOD: America votes. Join the Election Day conversation with #MyVote2016 https://t.co/BWuiwAxas6
ednewsdaily|educationviews|-0.4215|0.141|0.859|0.0|"PAC Tied to Teach for America Spends Big on a Local Indiana Election, but No One Quite https://t.co/jQ1sMzHedP https://t.co/c6YAh3RSgQ"
raincoaster|desertbunny|0.6418|0.0|0.654|0.346|RT @desertbunny: Newsrooms are so fun on election night
jesylroche|evanmcmurry|0.0|0.0|1.0|0.0|"RT @evanmcmurry: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
jesylroche||0.0|0.0|1.0|0.0|"RT @evanmcmurry: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
itsjustsadeen|Jena_Hammad|0.6369|0.0|0.682|0.318|@Jena_Hammad best thing to happen to you on election day
simxsimba_|isaatavares_|0.0|0.0|1.0|0.0|"RT @isaatavares_: putting it into spongebob terms, this is America before and after the election https://t.co/818HdJu06a"
simxsimba_|twitter|0.0|0.0|1.0|0.0|"RT @isaatavares_: putting it into spongebob terms, this is America before and after the election https://t.co/818HdJu06a"
bblancoynot|realDonaldTrump|0.0|0.0|1.0|0.0|"RT @realDonaldTrump: Before my FINAL campaign speech, I will get a list of Election Day Donors! Donate NOW! https://t.co/iZjo4q2gYA https:/"
bblancoynot|secure|0.0|0.0|1.0|0.0|"RT @realDonaldTrump: Before my FINAL campaign speech, I will get a list of Election Day Donors! Donate NOW! https://t.co/iZjo4q2gYA https:/"
maryzimnik|GuardianUS.|0.6369|0.0|0.792|0.208|Best place to get the #returns: @GuardianUS. Follow live #Election2016 updates as #votes come in | #ImWithHer    https://t.co/gJ2xFimRPK
maryzimnik|theguardian|0.6369|0.0|0.792|0.208|Best place to get the #returns: @GuardianUS. Follow live #Election2016 updates as #votes come in | #ImWithHer    https://t.co/gJ2xFimRPK
xDesiraee|smackingghoes|0.3818|0.129|0.588|0.282|RT @smackingghoes: either way we're all fcked no matter who wins the election
mlrandaaa|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
mlrandaaa|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
Erbibou|TheSimpsons|0.0|0.0|1.0|0.0|RT @TheSimpsons: ICYMI- Marge and Homer discuss the election. Watch! #TheSimpsonshttps://t.co/SwJP72VMft
DrBenWhitham|dmuleicester|0.0|0.0|1.0|0.0|RT @dmuleicester: #ElectionDay: DMU expert predicts the first 100 days for Trump &amp; Clinton: https://t.co/e8Zo6qWhYr https://t.co/2pRMHGA1kH
DrBenWhitham|dmu|0.0|0.0|1.0|0.0|RT @dmuleicester: #ElectionDay: DMU expert predicts the first 100 days for Trump &amp; Clinton: https://t.co/e8Zo6qWhYr https://t.co/2pRMHGA1kH
nerdfox|broadcast|0.0|0.0|1.0|0.0|Today's Elevate The Vote meditation for the 2016 election was deep. #ElevateTheVote  https://t.co/M04wqYfGF8
aNickel4thought|dyfl|0.0|0.0|1.0|0.0|"RT @dyfl: Just when you think this election cannot possibly offer up any more gifts to the meme economy, here comes Cake Trump"
JoSheram|jerome_corsi|-0.5859|0.153|0.847|0.0|RT @jerome_corsi: TRUMP NEEDS ALL POSSIBLE VOTERS IN PA - voter fraud being reported EVENING HOURS WILL DECIDE ELECTION - get all Trump vot
HollyWOhlweiler|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
decakarjeffrey|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
Blonde_Haleyyyy|G_Eazy|0.7644|0.0|0.752|0.248|"RT @G_Eazy: PLEASE GO OUT AND VOTE WHATEVER YOU DO, THIS COULD BE THE MOST IMPORTANT ELECTION OF OUR LIVES #imwithher #fuckdonaldtrump"
MichaelSticha1|Mozerik|0.0|0.0|1.0|0.0|RT @Mozerik: Election night starter kit https://t.co/t1tw2TXDGu
MichaelSticha1|twitter|0.0|0.0|1.0|0.0|RT @Mozerik: Election night starter kit https://t.co/t1tw2TXDGu
angieflyte99|keepingsanewth4|-0.2924|0.179|0.821|0.0|@keepingsanewth4 @jimsciutto It's not clear if it's election related...so there's that 
bryantre|TEDchris|0.0816|0.187|0.537|0.276|"RT @TEDchris: After this brutal election, can America heal? Psychologist @jonhaidt offered me some wisdom https://t.co/qN80oFDWcu Pls share!"
bryantre||0.0816|0.187|0.537|0.276|"RT @TEDchris: After this brutal election, can America heal? Psychologist @jonhaidt offered me some wisdom https://t.co/qN80oFDWcu Pls share!"
HannahHoelzen|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
BryanLarson3|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
BryanLarson3|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
FarmerGedon|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
FarmerGedon|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
natashafaith16|chasegoehring|0.5267|0.0|0.839|0.161|RT @chasegoehring: People are acting like this election is the end of the world ...We aren't getting nuked YET okay we still have some ti
Cheekie368|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
Cheekie368||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
MissLiberty1776|BoSnerdley|-0.4767|0.171|0.829|0.0|RT @BoSnerdley: WikiLeaks says it was under 'unrelenting' cyber attack on Election Day https://t.co/kf31Wxmlad via @MailOnline
MissLiberty1776|dailymail|-0.4767|0.171|0.829|0.0|RT @BoSnerdley: WikiLeaks says it was under 'unrelenting' cyber attack on Election Day https://t.co/kf31Wxmlad via @MailOnline
CohenBohen|Phil_Lewis_|0.5719|0.0|0.802|0.198|"RT @Phil_Lewis_: In a perfect world, this is how we would actually decide the election  #ElectionDay https://t.co/nnchd0Hymd"
CohenBohen|twitter|0.5719|0.0|0.802|0.198|"RT @Phil_Lewis_: In a perfect world, this is how we would actually decide the election  #ElectionDay https://t.co/nnchd0Hymd"
snowwhite_4|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Polls are closing in parts of nine states at 7 p.m. EST. Live results here: https://t.co/vLnb2jNCF6 https://t.co/a3fzaE
snowwhite_4|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Polls are closing in parts of nine states at 7 p.m. EST. Live results here: https://t.co/vLnb2jNCF6 https://t.co/a3fzaE
Dr_Straker|CNN's|-0.4767|0.341|0.659|0.0|I still only fucks with @CNN's Election coverage.
EnlightBystand|lizacsg|0.0|0.0|1.0|0.0|"RT @lizacsg: sometimes the election gets me down. but then, cheese. https://t.co/HG8AFl3igl"
EnlightBystand|twitter|0.0|0.0|1.0|0.0|"RT @lizacsg: sometimes the election gets me down. but then, cheese. https://t.co/HG8AFl3igl"
stringtheories|knitcollage|0.4199|0.0|0.763|0.237|I'm ready! Let the election coverage begin. @knitcollage @knitbaahpurl https://t.co/yaD9iRptAv
stringtheories|facebook|0.4199|0.0|0.763|0.237|I'm ready! Let the election coverage begin. @knitcollage @knitbaahpurl https://t.co/yaD9iRptAv
attheUC|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
Volla1Volland|CNNPolitics|0.0|0.0|1.0|0.0|RT @CNNPolitics: The first polls are closing at 7 p.m. ET. Get the latest results here https://t.co/jOauYyVeuX https://t.co/inPimatat2
Volla1Volland|cnn|0.0|0.0|1.0|0.0|RT @CNNPolitics: The first polls are closing at 7 p.m. ET. Get the latest results here https://t.co/jOauYyVeuX https://t.co/inPimatat2
NoshFoodandWine|nytimes|0.0|0.0|1.0|0.0|The Emotion of a Historic Vote https://t.co/pX0jiUMjCu
GrayDeenShaka|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
GrayDeenShaka|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
merinduh|latimes|0.0|0.0|1.0|0.0|@latimes shooting had nothing to do with election other than being near a local polling place. And it's AZUSA.
darf_69|IZOD|0.296|0.0|0.885|0.115|RT @IZOD: Share your voice this election. Make a statement with #MyVote2016 and Ken Bone in a red sweater. https://t.co/QX9fLqDpAL
darf_69|twitter|0.296|0.0|0.885|0.115|RT @IZOD: Share your voice this election. Make a statement with #MyVote2016 and Ken Bone in a red sweater. https://t.co/QX9fLqDpAL
fooIishshawn|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
fooIishshawn|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
thecattribe|MotherJones|0.0|0.0|1.0|0.0|RT @MotherJones: It's Election Day and Fox News Just Had a Total Meltdown https://t.co/NPdKw2zSHC https://t.co/lmawPdWCf9
thecattribe|motherjones|0.0|0.0|1.0|0.0|RT @MotherJones: It's Election Day and Fox News Just Had a Total Meltdown https://t.co/NPdKw2zSHC https://t.co/lmawPdWCf9
tkamins123|RealDJTrumpTeam|0.2124|0.0|0.934|0.066|"RT @RealDJTrumpTeam: Don't let up, get out to vote - this election is FAR FROM OVER! We are doing well but there is much time left. GO #FLO"
AlisshaM|LaurenJauregui|0.4795|0.0|0.881|0.119|RT @LaurenJauregui: I'm so excited that I was able to exercise my vote as a Cuban American Woman for the first time in this particular elec
DemsAbroad|amandamohar|0.0|0.0|1.0|0.0|RT @amandamohar: HK election watch location #1 checking in! @DemsAbroad #electionnight #ElectionNightAbroad https://t.co/kk6hPMG824
DemsAbroad|twitter|0.0|0.0|1.0|0.0|RT @amandamohar: HK election watch location #1 checking in! @DemsAbroad #electionnight #ElectionNightAbroad https://t.co/kk6hPMG824
mariizzle_|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
Mrlnzb|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
cupcake_queen97|dcexaminer|0.0|0.0|1.0|0.0|RT @dcexaminer: The first polls in Florida are about to close. Full state closings and our live electoral map: https://t.co/Iz2vhOwGcW #Ele
cupcake_queen97|washingtonexaminer|0.0|0.0|1.0|0.0|RT @dcexaminer: The first polls in Florida are about to close. Full state closings and our live electoral map: https://t.co/Iz2vhOwGcW #Ele
brianhoward41|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
tarintowers|edbott|-0.7964|0.372|0.628|0.0|@edbott my biggest fear about this election is that someone would die of it.
kara_klimekk|RealHeatherRoss|0.0|0.0|1.0|0.0|RT @RealHeatherRoss: When you're two weeks away from rigging an election and then the FBI reopens your investigation. https://t.co/w0GMEHG0
kara_klimekk|t|0.0|0.0|1.0|0.0|RT @RealHeatherRoss: When you're two weeks away from rigging an election and then the FBI reopens your investigation. https://t.co/w0GMEHG0
3beansalad|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
_baileefox_|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
_baileefox_|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
megasafeinvest|reuters|0.0|0.0|1.0|0.0|"Stocks, Mexican peso climb ahead of US election results - Reuters https://t.co/qNEyNfxkFQ"
ONLYTRUMP4USA|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
blackwood_julie|DavidCornDC|-0.7096|0.312|0.688|0.0|RT @DavidCornDC: I have been banned by @realDonaldTrump. I was denied credentials for Trump election night event.
ackwdw123|it|0.0|0.0|1.0|0.0|4chan May Have Brought Down Pro-Clinton Phone Lines Before Election Day https://t.co/BkLpuZxOx2
Shelbscarps|Gizmodo|0.0|0.0|1.0|0.0|RT @Gizmodo: The polls close in six states in just 15 minutes. Here's how to watch the Election Night returns streaming live https://t.co/S
Shelbscarps|jack|0.0|0.0|1.0|0.0|RT @Gizmodo: The polls close in six states in just 15 minutes. Here's how to watch the Election Night returns streaming live https://t.co/S
ScottFralick|JHertnerCTV|0.0|0.0|1.0|0.0|RT @JHertnerCTV: Nap  .. time for some edge of the seat election watching #ElectionParty #Merica #RealLifeRealityShow #NewEra
mlogika1|abcnews|0.25|0.0|0.867|0.133|RT @abcnews: .@HillaryClinton one step away from snaring her dream job #Election2016 https://t.co/XpMh9z93OP https://t.co/mPAFkHucrD
mlogika1|abc|0.25|0.0|0.867|0.133|RT @abcnews: .@HillaryClinton one step away from snaring her dream job #Election2016 https://t.co/XpMh9z93OP https://t.co/mPAFkHucrD
ProLivid|twitter|0.0|0.0|1.0|0.0|This year's election  https://t.co/pAVGg2kLH7
thesaadahmed|LBC|0.0|0.0|1.0|0.0|"RT @LBC: .@ChukaUmunna tells Iain he's hearing tonight from people involved in the US election ""it's very tight"" https://t.co/4zu41YcSJD ht"
thesaadahmed|lbc|0.0|0.0|1.0|0.0|"RT @LBC: .@ChukaUmunna tells Iain he's hearing tonight from people involved in the US election ""it's very tight"" https://t.co/4zu41YcSJD ht"
Twisty58|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
USAncestors1636|POTUS|0.5709|0.0|0.802|0.198|@POTUS  Barack Obama is now viewed more positively than Ronald Reagan was in 1988 #election  https://t.co/JhITpM6uiJ
USAncestors1636|washingtonpost|0.5709|0.0|0.802|0.198|@POTUS  Barack Obama is now viewed more positively than Ronald Reagan was in 1988 #election  https://t.co/JhITpM6uiJ
smallant|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
smallant|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
TLVRP_Tennessee|wjhl|0.0|0.0|1.0|0.0|"#Tennessee #Memphis #Nashville LIVE UPDATES: November 8 local, state election results https://t.co/D0p3cq09t9"
AshleyyOwnby|TweetLikeAGirI|0.6249|0.0|0.661|0.339|RT @TweetLikeAGirI: A great way to start Election Day https://t.co/RpgZgjX3lG
AshleyyOwnby|twitter|0.6249|0.0|0.661|0.339|RT @TweetLikeAGirI: A great way to start Election Day https://t.co/RpgZgjX3lG
alenaangel16|raaaqcity|0.5707|0.0|0.817|0.183|"RT @raaaqcity: please exercise your right to vote tomorrow! unless you're a trump supporter, then election day is on nov. 28th for you guys"
JR818FL|abcnews|0.0|0.0|1.0|0.0|2016 Presidential Election Results: Live Map - ABC News https://t.co/TxHjYY39VV
h8breeding|CherOfficiaI|0.6633|0.0|0.783|0.217|RT @CherOfficiaI: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
oxnfre|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
juliarosexox|Powerful|0.7085|0.0|0.734|0.266|"RT @Powerful: Me @ the beginning of the election: Ain't no way America letting a cheeto become president. lol what a joke Me November 8,"
wmarsburg|mrchrisaddison|-0.4118|0.116|0.884|0.0|"RT @mrchrisaddison: The last time I was watching a US election this tense, I was standing in the room with Selina Meyer and her team."
zauxier|jimgeraghty|0.7351|0.0|0.714|0.286|"RT @jimgeraghty: The Trump party victory cake. This election is like a surreal, twisted dream where nothing makes sense and its taking f"
qamaranissa|chefalexander1|0.0|0.0|1.0|0.0|"RT @chefalexander1: If I could vote this election, I would. #ImWithHer"
NoYardstick|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
NoYardstick|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
Sebai2s|cnnpolitics|0.0|0.0|1.0|0.0|"CNN: 2016 presidential election, House, Senate results via @cnnpolitics https://t.co/DZXRbM2lx8"
Sebai2s|edition|0.0|0.0|1.0|0.0|"CNN: 2016 presidential election, House, Senate results via @cnnpolitics https://t.co/DZXRbM2lx8"
PatriciaFritz4|MotherJones|0.0|0.0|1.0|0.0|RT @MotherJones: It's Election Day and Fox News Just Had a Total Meltdown https://t.co/NPdKw2zSHC https://t.co/lmawPdWCf9
PatriciaFritz4|motherjones|0.0|0.0|1.0|0.0|RT @MotherJones: It's Election Day and Fox News Just Had a Total Meltdown https://t.co/NPdKw2zSHC https://t.co/lmawPdWCf9
jdbfttori|harIeystorm|-0.9199|0.346|0.591|0.062|"RT @harIeystorm: BERNIE JUST WANTED TO HELP, BUT YALL HAD TO LET THE CRIMINAL AND THE RACIST GO THROUGH TO THE ELECTION  #ElectionNight htt"
AliasHandler|MargHartmann|0.357|0.0|0.858|0.142|RT @MargHartmann: As if I werent jealous enough that my polling place doesnt do I voted stickers https://t.co/Kf8XoPXTpG
AliasHandler|vox|0.357|0.0|0.858|0.142|RT @MargHartmann: As if I werent jealous enough that my polling place doesnt do I voted stickers https://t.co/Kf8XoPXTpG
millie_heyyy|Markgatiss|-0.7096|0.362|0.467|0.171|"RT @Markgatiss: I have a dreadful, sick feeling of foreboding about the US election. I hope to Christ I'm wrong."
joabbess|nataliemjb|-0.8016|0.286|0.714|0.0|"RT @nataliemjb: So after all the hell of the last year, having a very boring election night would be very 2016."
justdolanit|EthanDolan|0.4572|0.0|0.864|0.136|@EthanDolan @GraysonDolan so curious to know this; who would you have voted for in the election if you could? #USElection2016
LyellBan|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
LyellBan|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
jhseher|CNNPolitics|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
jhseher|twitter|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
PhilDeCarolis|business|0.0|0.0|1.0|0.0|RT @business: We're live-blogging #ElectionNight. Follow along here as the results roll in https://t.co/HYCnbzTiqS https://t.co/D20AtkGCw6
PhilDeCarolis|bloomberg|0.0|0.0|1.0|0.0|RT @business: We're live-blogging #ElectionNight. Follow along here as the results roll in https://t.co/HYCnbzTiqS https://t.co/D20AtkGCw6
SculptNewYork|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
SculptNewYork||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
midnightdrivinn|godnhs|0.5023|0.0|0.84|0.16|"RT @godnhs: I know the election has everyone's attention, but I'd just like to remind you about this: https://t.co/8dB2eweFxO"
midnightdrivinn|twitter|0.5023|0.0|0.84|0.16|"RT @godnhs: I know the election has everyone's attention, but I'd just like to remind you about this: https://t.co/8dB2eweFxO"
outerspes|CALUMDATING|0.1571|0.115|0.737|0.147|RT @CALUMDATING: bless calum for tweeting about the election/voting even though he's not American + on holidays
roofusfirefly|ACLUaz|0.6833|0.0|0.789|0.211|"RT @ACLUaz: HUGE DEAL: If You Voted Early, Check to make sure it counted! 7k ballots in Maricopa Co. have issue https://t.co/VPmYTTyUWC via"
roofusfirefly|azcentral|0.6833|0.0|0.789|0.211|"RT @ACLUaz: HUGE DEAL: If You Voted Early, Check to make sure it counted! 7k ballots in Maricopa Co. have issue https://t.co/VPmYTTyUWC via"
joelwatts|instagram|0.4019|0.0|0.69|0.31|"Election Party Snacks: Republican Raspberries, Democratic https://t.co/RFekpJBDv2"
Radhika0Sharma|itsHIMYMquotes|0.0|0.0|1.0|0.0|RT @itsHIMYMquotes: Since it's Election Day... https://t.co/IEFE9jhYVT
Radhika0Sharma|twitter|0.0|0.0|1.0|0.0|RT @itsHIMYMquotes: Since it's Election Day... https://t.co/IEFE9jhYVT
tillymomma21|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
ekimballin|GabMeoww|0.3612|0.0|0.902|0.098|RT @GabMeoww: This election is like waiting for Christmas morning... You could get a lump of coal or grandma gives you the same sweater as
sjwjs|billmckibben|0.4404|0.0|0.873|0.127|RT @billmckibben: New numbers just in: 93% of the good things about this election had to do with that guy @BernieSanders
iStigrrr|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
boisvert813|untappd!|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/ioF5fKjThm #voteforbeer
boisvert813|untappd|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/ioF5fKjThm #voteforbeer
Goodyear29|penguins|0.2716|0.0|0.793|0.207|@penguins game is more important than this election bs
TLVRP_Tennessee|oakridger|0.1027|0.117|0.748|0.136|#Tennessee #Memphis #Nashville Trump spent a good portion of Election Day sowing doubt about the legitimacy of the https://t.co/fy868izwPk
madisonjheath_|garyfromteenmom|0.7579|0.0|0.683|0.317|RT @garyfromteenmom: there should be a gender reveal party instead of announcing the winner of the election
billionairesson|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
MizCoretta|RedApplePol|0.5473|0.0|0.531|0.469|RT @RedApplePol: HERE'S HOPING  https://t.co/v0Yvnpt9hh
MizCoretta|aljazeera|0.5473|0.0|0.531|0.469|RT @RedApplePol: HERE'S HOPING  https://t.co/v0Yvnpt9hh
FightNightatJoe|ahtrapsm|0.2732|0.0|0.884|0.116|@ahtrapsm to try as well. We're covering this about as heavily as if it was a Norwegian election
BuzzFeed|buzzfeed|0.6115|0.0|0.734|0.266|People are stress-eating the most delicious treats before the election https://t.co/6p2zZ7oVdg https://t.co/eVl1SfBk7B
SternishOwl|curtisstigers|-0.7798|0.254|0.746|0.0|RT @curtisstigers: Hey @mrjamesob I just found this wanker creeping around our election &amp; mumbling nonsense. Does he belong to you guys? ht
EEGRC98|0hour|0.0|0.0|1.0|0.0|RT @0hour: https://t.co/2S72Q1xk2DIndiana70% as of nowits happening!
EEGRC98|t|0.0|0.0|1.0|0.0|RT @0hour: https://t.co/2S72Q1xk2DIndiana70% as of nowits happening!
DeeDeeMarberry|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
Castaneda1210|Capitals|0.0|0.0|1.0|0.0|Im Tweeting to #VoteHoltby for @Capitals bobblehead night! Visit https://t.co/I595bu6URX for more details! #CapsElectionNight
Castaneda1210|nhl|0.0|0.0|1.0|0.0|Im Tweeting to #VoteHoltby for @Capitals bobblehead night! Visit https://t.co/I595bu6URX for more details! #CapsElectionNight
kmcmahon44|barstoolsports|0.5719|0.0|0.856|0.144|"RT @barstoolsports: Before you move to Canada after this election, learn some more about our neighbors to the north. They're happy to have"
scoj24|YahooSports|0.0|0.0|1.0|0.0|RT @YahooSports: Ric Flair voted for exactly who you'd think Ric Flair would vote for: Ric Flair. https://t.co/2GceP31bit https://t.co/wI6G
scoj24|sports|0.0|0.0|1.0|0.0|RT @YahooSports: Ric Flair voted for exactly who you'd think Ric Flair would vote for: Ric Flair. https://t.co/2GceP31bit https://t.co/wI6G
Pinkychelle|YouTube|-0.5962|0.297|0.578|0.125|"I liked a @YouTube video from @weallbe https://t.co/GmUfxDbQVJ ""Baba Dick GREgory: THE GaME's BEen Rigged!!! Election Eve 2016"
Pinkychelle|youtube|-0.5962|0.297|0.578|0.125|"I liked a @YouTube video from @weallbe https://t.co/GmUfxDbQVJ ""Baba Dick GREgory: THE GaME's BEen Rigged!!! Election Eve 2016"
SimplyyRosee|AnimeUproar|0.0|0.0|1.0|0.0|RT @AnimeUproar: We are going LIVE - Election 2016 (ANIME EDITION) -  https://t.co/7cXkLGIyuy #anime #ElectionDay #ElectionNight #Elections
SimplyyRosee|youtube|0.0|0.0|1.0|0.0|RT @AnimeUproar: We are going LIVE - Election 2016 (ANIME EDITION) -  https://t.co/7cXkLGIyuy #anime #ElectionDay #ElectionNight #Elections
ginnyv58|TheMarkRomano|0.0516|0.102|0.789|0.109|RT @TheMarkRomano: It is a real problem that so much rides on one Presidential election.It should not be this way.We are truly at the p
paulrlanni|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Deplorablecasee|DonaldJTrumpJr|0.3164|0.0|0.906|0.094|RT @DonaldJTrumpJr: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERSGET OUT AND VOTE! Find 5 others. This is our chance to take back Am
Unlaiga|NextGenPhoenix|-0.5423|0.132|0.868|0.0|RT @NextGenPhoenix: This Election brought out the bad in my city. Places got shut down by mass shootings. First time taking bullets for unp
TheUndine3|10thAmendment|-0.7342|0.262|0.668|0.07|@10thAmendment @angelinthepine psyop false flag. Government will do anything even kill us to rig election. Vote!!! Don't let them stop you
NadineORegan|MsAmyHerron|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
NadineORegan|theguardian|0.0|0.0|1.0|0.0|RT @MsAmyHerron: The only link you need right now https://t.co/HnGEb3QhNk #ElectionNight
Gig74Hgig|maramcewin|0.0|0.0|1.0|0.0|RT @maramcewin: Daughter just made our election signs for tonight's election party#ElectionNight #Election2016 #nyvotes @HillaryCl
realtor99587|realtor101blog|0.6052|0.0|0.767|0.233|Election? What Election?! Check Out These Cute Animals We Found in ListingPhotos! https://t.co/O7hFdfbhjv https://t.co/WUHglMwmNb
fortymileFrank|fernacarieles|0.6523|0.1|0.651|0.249|"RT @fernacarieles: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://"
fortymileFrank||0.6523|0.1|0.651|0.249|"RT @fernacarieles: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://"
greenlawley|lovelaurenxjenn|0.5719|0.0|0.821|0.179|RT @lovelaurenxjenn: If Trump or Hillary  Wins The Election I Am Moving  Out Of The Country  Goodbye America  Hello   N
krystalstory|Cronkite_ASU|0.0|0.0|1.0|0.0|RT @Cronkite_ASU: Walter Cronkite on election night. #CronkiteAt100 https://t.co/pqzgddeELd
krystalstory|twitter|0.0|0.0|1.0|0.0|RT @Cronkite_ASU: Walter Cronkite on election night. #CronkiteAt100 https://t.co/pqzgddeELd
mayadiez|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
PASSMAN47|charliekirk11|0.1779|0.108|0.757|0.135|RT @charliekirk11: To my fellow millennials: don't vote for someone who will enrich herself &amp; gain political power - reject career politici
FloMOUVAUX|Jonbuckhouse|0.6239|0.0|0.843|0.157|RT @Jonbuckhouse: The Polls are starting to close all over the US! Who do you think will win the election?  #ElectionNight #electionday #iV
libbytubbergen|WMUSocial|-0.6229|0.29|0.71|0.0|RT @WMUSocial: Fuck the election! Broncos about to go 10-r0w tonight!
EJRifkind|Yair_Rosenberg|0.5719|0.0|0.778|0.222|"RT @Yair_Rosenberg: Whatever else has happened this election, I am thankful for this moment. https://t.co/guDLhsRptO"
EJRifkind|twitter|0.5719|0.0|0.778|0.222|"RT @Yair_Rosenberg: Whatever else has happened this election, I am thankful for this moment. https://t.co/guDLhsRptO"
casheyesblond|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
casheyesblond|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
NancyIncocoa|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
webcentraltv|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
webcentraltv|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
JWarren5180|Franklin_Graham|0.765|0.0|0.714|0.286|RT @Franklin_Graham: This election isnt overits going to be a tight race. Join with family or friends to pray throughout the night that
esmerugh|CherOfficiaI|0.6633|0.0|0.783|0.217|RT @CherOfficiaI: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
jalenalizabeth|whats_up_Erv|0.3612|0.0|0.884|0.116|"RT @whats_up_Erv: Thank the lord for women voting sticker selfies on Instagram, never would have known today was the election."
jenny_rusher22|KeeganAllen|0.6249|0.0|0.843|0.157|"RT @KeeganAllen: Instead of looking at this election as a series finale of the Great American reality show, look at it as your life...start"
RhondellaW|WDFx2EU8|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
RhondellaW|t|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
zakcreative|TheDailyShow|0.0|0.0|1.0|0.0|RT @TheDailyShow: Election Day is here. Get out and vote. https://t.co/C5rqe8KTyt https://t.co/BKHBkUjtn7
zakcreative|cc|0.0|0.0|1.0|0.0|RT @TheDailyShow: Election Day is here. Get out and vote. https://t.co/C5rqe8KTyt https://t.co/BKHBkUjtn7
leftcobain|skilletmusic|-0.3595|0.122|0.878|0.0|RT @skilletmusic: Skillet is the 1st Christian band to hit No. 1 on the Mainstream Rock Chart with #FeelInvincible! https://t.co/acdfzlImhg
leftcobain|skillet|-0.3595|0.122|0.878|0.0|RT @skilletmusic: Skillet is the 1st Christian band to hit No. 1 on the Mainstream Rock Chart with #FeelInvincible! https://t.co/acdfzlImhg
EceeR___|ImageSlays|-0.1531|0.096|0.904|0.0|RT @ImageSlays: If Donald Trump Looses the election I'll give everybody who RTs this $5 PayPal.
PHES_ITC|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
PHES_ITC|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
Pas_Normal|TBNSport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
Pas_Normal|tbnsport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
AngelNapoles4|DonaldJTrumpJr|0.69|0.0|0.802|0.198|RT @DonaldJTrumpJr: Friends sending me pics and lots of calls about long lines. Please wait it out and VOTE! Every vote is needed. Your VOI
JimbauxsJournal|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
JimbauxsJournal|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
WandaAlbright1|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: Kai sporting the #MAGA hat. She has only asked 300 times today if she could go vote. Not yet! But YOU CAN! Go Vote!!! #
PaceTire|RollTribe2016|-0.6249|0.339|0.661|0.0|@RollTribe2016 this election brought out the worst in people
RoneyCarias|YouTube|0.4215|0.0|0.811|0.189|I liked a @YouTube video from @theyoungturks https://t.co/icFeAIzwF5 The Young Turks Election Day Coverage 2016
RoneyCarias|youtube|0.4215|0.0|0.811|0.189|I liked a @YouTube video from @theyoungturks https://t.co/icFeAIzwF5 The Young Turks Election Day Coverage 2016
tatumdeems|KilgoreMicah|0.6597|0.0|0.803|0.197|"RT @KilgoreMicah: Christians, we're already free in the Lord. whatever the outcome of this election may be, rest in the fact that God reign"
Tolu__A|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Tolu__A|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
biebertopping|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
biebertopping|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
NickDawybida|missmazzz|0.0|0.0|1.0|0.0|RT @missmazzz: I just voted!!! In the presidential election!!! I'm a real life grownup!!!
jwilson195506|NBCNewsPR|-0.4019|0.144|0.856|0.0|RT @NBCNewsPR: BOOKMARK: @NBCNews Battleground Map https://t.co/YAWPTcaBqvTune in to #Decision2016 tonight on @NBC beginning at 7p ET #
jwilson195506|t|-0.4019|0.144|0.856|0.0|RT @NBCNewsPR: BOOKMARK: @NBCNews Battleground Map https://t.co/YAWPTcaBqvTune in to #Decision2016 tonight on @NBC beginning at 7p ET #
vasquez_sari|Dan_Juarez_|0.4939|0.0|0.714|0.286|RT @Dan_Juarez_: In honor of the election today https://t.co/EKStC0TGcU
vasquez_sari|twitter|0.4939|0.0|0.714|0.286|RT @Dan_Juarez_: In honor of the election today https://t.co/EKStC0TGcU
PepeAnabolic|Fash_UK|0.2716|0.0|0.861|0.139|RT @Fash_UK: Imagine not voting in the most important election of our lifetime.... WEW
JadeFrdrik|_Gorran|0.0|0.0|1.0|0.0|"RT @_Gorran: This election affects all of us, and so many people don't seem to understand. #ElectionDay"
chicken_nuggit|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
chicken_nuggit|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
PaulMakesMovies|TIME|0.4019|0.0|0.856|0.144|RT @TIME: Mixed Drinks are $13 and beer is $11 at Donald Trump's election night party https://t.co/GqEEQDeBCf
PaulMakesMovies|fortune|0.4019|0.0|0.856|0.144|RT @TIME: Mixed Drinks are $13 and beer is $11 at Donald Trump's election night party https://t.co/GqEEQDeBCf
irasroom|nytimes|0.0|0.0|1.0|0.0|"RT @nytimes: Live 2016 election results, as they come in https://t.co/Kir4tzdGWF https://t.co/ejeePNRkvG"
irasroom|nytimes|0.0|0.0|1.0|0.0|"RT @nytimes: Live 2016 election results, as they come in https://t.co/Kir4tzdGWF https://t.co/ejeePNRkvG"
dc3246|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
JmitchJon|realtor|0.6052|0.0|0.78|0.22|Election? What Election?! Check Out These Cute Animals We Found in Listing Photos! https://t.co/DgocnH9x4j https://t.co/reAZ5zy5wE
rafoleiro|theverge|0.0|0.0|1.0|0.0|10 provocative political novels to read after the election https://t.co/ugp6Zsjk8I
yin_naya|AmazingDanny_|0.5859|0.0|0.858|0.142|"RT @AmazingDanny_: Americans are yet to know the winner of today's election. If it was Nigeria, we for dun know the result before evening."
MrFijiWiji|JackBrommel|0.0|0.0|1.0|0.0|RT @JackBrommel: Reppin the obvious choice for this election  https://t.co/2L2fBdN3zU
MrFijiWiji|twitter|0.0|0.0|1.0|0.0|RT @JackBrommel: Reppin the obvious choice for this election  https://t.co/2L2fBdN3zU
usconsulatekhi|shareamerica|0.3595|0.0|0.889|0.111|RT @shareamerica: LIVE NOW: Election Night webchat w/ political experts answering ?s about the U.S. election process. Join the chat! https
justjaney_|nedfulmer|0.3182|0.0|0.859|0.141|"RT @nedfulmer: ""I just spellchecked election 5 times to make sure I didn't write erection"" -- @korndiddy"
tooshort__|drmoore|0.7845|0.0|0.717|0.283|"RT @drmoore: Well, it's almost over. What we can all agree on: anyone who has enjoyed this election year needs to seek counseling."
schmemmm|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
schmemmm|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
gocoo|LaurenJauregui|0.4795|0.0|0.881|0.119|RT @LaurenJauregui: I'm so excited that I was able to exercise my vote as a Cuban American Woman for the first time in this particular elec
mooovingmoments|live|0.0|0.0|1.0|0.0|Election 2016 https://t.co/NWnnL4ouMl
PhineasZest|Talkmaster|-0.5423|0.155|0.774|0.071|RT @Talkmaster: Election may be decided by voters who fled Democrat New England to GOP states and then voted to create the same hell they f
marioterrones25|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
marioterrones25|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
stephgue7|Things4WhitePpl|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
stephgue7|twitter|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
GalipDalay|SharqForum|0.0|0.0|1.0|0.0|RT @SharqForum: What Does the U.S. Election Mean for the Middle East?https://t.co/xpC8PVCl55 https://t.co/6vyDRWsTNq
GalipDalay|sharqforum|0.0|0.0|1.0|0.0|RT @SharqForum: What Does the U.S. Election Mean for the Middle East?https://t.co/xpC8PVCl55 https://t.co/6vyDRWsTNq
yagirlcdollas|sariuhhh|0.4019|0.151|0.576|0.273|RT @sariuhhh: wow i'm like...genuinely nervous for these election results
MaryEBarnes|DRUDGE_REPORT|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
MaryEBarnes|businessinsider|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
DevloPM|SoaRPraizist|0.5719|0.0|0.802|0.198|"RT @SoaRPraizist: If Trump wins the election, I will make artwork for everyone that RTs this tweet"
Becky_LoveDemi|MichelleKrys|-0.7206|0.208|0.741|0.051|"RT @MichelleKrys: If you want something to keep your mind off the election, DEAD GIRLS SOCIETY is out today! https://t.co/bSAPWXBSVR https:"
Becky_LoveDemi|amazon|-0.7206|0.208|0.741|0.051|"RT @MichelleKrys: If you want something to keep your mind off the election, DEAD GIRLS SOCIETY is out today! https://t.co/bSAPWXBSVR https:"
Redheadedbird|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
EmmaHam2|allienolann|0.2732|0.0|0.92|0.08|RT @allienolann: just wanted to remind everyone that God already knows the outcome of the election &amp; that He is in control of His kingdom n
basedruba|dj_rocklee|0.5374|0.082|0.752|0.166|RT @dj_rocklee: Shiiitttt if Donald Trump wins this election im warning ALL YALL !!!!! Knuck if you buck white America. Knuck if you the
papiwhitelion|papiwhitelion|0.5719|0.0|0.812|0.188|RT @papiwhitelion: Will Bill Clinton be the 'First Man' of the USA if Hillary wins this Election?
CynthiaMace1|RMSilverman|0.0|0.0|1.0|0.0|RT @RMSilverman: FSN LIVE and TV Azteca reporting from NYC on the eve of the presidential election @FSNLIVE  @Azteca  @featurestory https:/
CynthiaMace1||0.0|0.0|1.0|0.0|RT @RMSilverman: FSN LIVE and TV Azteca reporting from NYC on the eve of the presidential election @FSNLIVE  @Azteca  @featurestory https:/
DOLORESVESTRICH|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
DOLORESVESTRICH|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
tevinclarke252|YouTube|0.0|0.0|1.0|0.0|The Young Turks Election Day Coverage 2016 https://t.co/F5xwQLGrYq via @YouTube
tevinclarke252|youtube|0.0|0.0|1.0|0.0|The Young Turks Election Day Coverage 2016 https://t.co/F5xwQLGrYq via @YouTube
JanLeeEmmer|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
thebizofmisery|ephrata|-0.2732|0.116|0.884|0.0|RT @ephrata: Just gonna drop this here so you can weigh your options on Election Day  https://t.co/vLImlUcvtU
thebizofmisery|twitter|-0.2732|0.116|0.884|0.0|RT @ephrata: Just gonna drop this here so you can weigh your options on Election Day  https://t.co/vLImlUcvtU
fordstokes|KarlRove|-0.4767|0.307|0.693|0.0|@KarlRove Unfair shot at Trump on Election night.
___jomeeee|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
TheSteveHolland|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
TheSteveHolland||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
aspen1031|blvckpapii|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
aspen1031|twitter|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
Restrepojuanfe|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
Restrepojuanfe|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
elmorephd|NRO|0.0|0.0|1.0|0.0|"RT @NRO: Early Exit Polls: Trump Opens YUGE Gap between College-Educated, Non-College-Educated Whiteshttps://t.co/ADpCNhYfiC #ElectionNight"
djrobdipaolo|instagram|-0.2547|0.197|0.7|0.103|"Ok Presidential Election, I don't like you and you don't like me. Let's just get through this so https://t.co/6VTJHFB2Jf"
drew4524|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
nwi_kerrye|instagram|-0.4973|0.297|0.703|0.0|There's nothing like Election Night pizza in the newsroom. It's like https://t.co/2HRCnoqwQ0
babiplant|petesmoonbase|-0.2466|0.193|0.664|0.143|RT @petesmoonbase: Feels more like a bad reality tv show than an actual presidential election  #ElectionNight
kimgee41|joshmancuso|0.0|0.0|1.0|0.0|RT @joshmancuso: Today I voted for @Evan_McMullin. It's a vote for conservative principles and for our future. #Election
kirstenp998|kurtsteiss|0.0|0.0|1.0|0.0|"RT @kurtsteiss: There are now 6,884 flags on the #okstate library lawn, and they aren't for the election. Each flag represents a soldier ki"
wtfstavo|LaurenJauregui|0.4795|0.0|0.881|0.119|RT @LaurenJauregui: I'm so excited that I was able to exercise my vote as a Cuban American Woman for the first time in this particular elec
MWatsPatriot|nbcconnecticut|0.0|0.0|1.0|0.0|#trumpI just told #NBCCT I voted today for Donald #Trump. Follow @nbcconnecticut for the latest election news. https://t.co/IX8mb1stcJ
MWatsPatriot|nbcconnecticut|0.0|0.0|1.0|0.0|#trumpI just told #NBCCT I voted today for Donald #Trump. Follow @nbcconnecticut for the latest election news. https://t.co/IX8mb1stcJ
sisterbarbieq|marinanachos|0.4939|0.0|0.802|0.198|RT @marinanachos: How early is too early for Election Day drinking?  Asking for a friend.
MarboGarbo|HIGH_TIMES_Mag|0.2225|0.0|0.921|0.079|RT @HIGH_TIMES_Mag: We're back on FB Live! Want to know the second weed gets legalized? IGH TIMES is covering the election live! https://t.
MarboGarbo||0.2225|0.0|0.921|0.079|RT @HIGH_TIMES_Mag: We're back on FB Live! Want to know the second weed gets legalized? IGH TIMES is covering the election live! https://t.
xlovelyfranta|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
xlovelyfranta|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
gpena|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
Synbane|tylissius|-0.3382|0.298|0.527|0.176|"@tylissius Jokes on you, the election fucks you!"
NotChrisWells|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
neatIester|StanceFrac|0.5719|0.0|0.791|0.209|RT @StanceFrac: If Donald trump wins the election I'll PayPal everyone that rted this $1
yourbeth_friend|TamEdwards6abc|0.4939|0.0|0.862|0.138|"RT @TamEdwards6abc: Women are flocking to Susan B Anthony's NY State gravesite, leaving their ""I Voted"" stickers on headstone, in honor of"
SOgnenis|ElementsMatter|0.0|0.0|1.0|0.0|RT @ElementsMatter: 2016 Election Night: Live coverage and results | FiveThirtyEight https://t.co/JkhpQqLMUr
SOgnenis|fivethirtyeight|0.0|0.0|1.0|0.0|RT @ElementsMatter: 2016 Election Night: Live coverage and results | FiveThirtyEight https://t.co/JkhpQqLMUr
BorisNotDJ|jermainenyc|0.5936|0.0|0.805|0.195|"can't wait till this election is over..So we can talk about more important things, like my bday bash w/@jermainenyc this Fri @schimanskinyc"
DJ_Homewrecker|DJ_Homewrecker|-0.5319|0.209|0.791|0.0|RT @DJ_Homewrecker: TRUMP IS ABOUT TO LOSE AN ELECTION ON TACO TUESDAY. SO FITTING.
zengirl55|ananavarro|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
zengirl55|twitter|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
IdeaGov|jacobsoboroff|0.3182|0.0|0.892|0.108|RT @jacobsoboroff: Huge lines at this Philly polling place with less than two hours to go until polls close.  https://t.co/nrQfFAMk1Q
IdeaGov|twitter|0.3182|0.0|0.892|0.108|RT @jacobsoboroff: Huge lines at this Philly polling place with less than two hours to go until polls close.  https://t.co/nrQfFAMk1Q
KoolaidUSA|NewYorker|0.4588|0.0|0.842|0.158|RT @NewYorker: The Trump campaign was laughed out of the courtroom in Nevada today. https://t.co/XpavP0b3k8 #ElectionDay https://t.co/hmjmK
KoolaidUSA|newyorker|0.4588|0.0|0.842|0.158|RT @NewYorker: The Trump campaign was laughed out of the courtroom in Nevada today. https://t.co/XpavP0b3k8 #ElectionDay https://t.co/hmjmK
StellaLelohan|BreitbartNews|0.802|0.0|0.631|0.369|"Reuters Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader'  https://t.co/oQwv6k1xu9 via @BreitbartNews"
StellaLelohan|breitbart|0.802|0.0|0.631|0.369|"Reuters Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader'  https://t.co/oQwv6k1xu9 via @BreitbartNews"
djajiprime|squalloogal|0.0|0.0|1.0|0.0|RT @squalloogal: Only place to get the facts on this election and what's to come #tytlive https://t.co/2phE3aPrCi
djajiprime|twitter|0.0|0.0|1.0|0.0|RT @squalloogal: Only place to get the facts on this election and what's to come #tytlive https://t.co/2phE3aPrCi
ranpaq|HalleyBorderCol|0.7703|0.0|0.74|0.26|"RT @HalleyBorderCol: For anyone wanting election results as them come in, the Guardian site seems quite good. Looking good for #Trump!htt"
mae_claire1|GAVlNREACTS|0.6249|0.0|0.661|0.339|RT @GAVlNREACTS: A great way to start Election Day https://t.co/yr6QAP3orF
mae_claire1|twitter|0.6249|0.0|0.661|0.339|RT @GAVlNREACTS: A great way to start Election Day https://t.co/yr6QAP3orF
NC1Sam|NewsCenter1|-0.5423|0.189|0.723|0.088|Poll workers say it's been a smooth day at Pinedale Elementary for voters. Join us on @NewsCenter1 for tonight's fu https://t.co/VqLSTOqV89
NC1Sam|twitter|-0.5423|0.189|0.723|0.088|Poll workers say it's been a smooth day at Pinedale Elementary for voters. Join us on @NewsCenter1 for tonight's fu https://t.co/VqLSTOqV89
MasonHartzell14|ColtonRamos|0.3818|0.0|0.822|0.178|RT @ColtonRamos: The only man who can protect us from this election  https://t.co/U7A0c5Oa6P
MasonHartzell14|twitter|0.3818|0.0|0.822|0.178|RT @ColtonRamos: The only man who can protect us from this election  https://t.co/U7A0c5Oa6P
ObjectiviTweets|ariarmstrong|0.4404|0.0|0.805|0.195|"RT @ariarmstrong: 538 has a good live blog going of the election, btw: https://t.co/dxzoPHZiZk"
ObjectiviTweets|fivethirtyeight|0.4404|0.0|0.805|0.195|"RT @ariarmstrong: 538 has a good live blog going of the election, btw: https://t.co/dxzoPHZiZk"
koalagirl08|dressed_sharp|-0.7707|0.324|0.676|0.0|"RT @dressed_sharp: There s nothing patriotic about accepting a fraudulent election, real Americans will go to court if #trump loses because"
EffortlessChick|twitter|-0.5106|0.32|0.68|0.0|I'm sick of it... Election go away https://t.co/Jw5Uc3KoXE
elaineprettyeye|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
honeynutlexios|InappropriateSB|0.0|0.0|1.0|0.0|RT @InappropriateSB: This election in a nutshell https://t.co/TE1m8Scmmi
honeynutlexios|twitter|0.0|0.0|1.0|0.0|RT @InappropriateSB: This election in a nutshell https://t.co/TE1m8Scmmi
Electric41E|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: WikiLeaks editor Julian Assange's statement today on the US election https://t.co/Q6KEChqm1B https://t.co/ZdZlolZJMl
Electric41E|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: WikiLeaks editor Julian Assange's statement today on the US election https://t.co/Q6KEChqm1B https://t.co/ZdZlolZJMl
El_Ma3stro77|lp_1516|0.0775|0.079|0.791|0.13|@lp_1516 @IZOD I didn't vote you know that lol cause I know it's important to do it but I don't think it's worth in this election
Ultimate_Solo|CNN|-0.1531|0.071|0.929|0.0|RT @CNN: Time is running out for @HillaryClinton &amp; @realDonaldTrump. Its a close race. Dont miss a moment on election night with CNN. htt
efairhurst|nbcphiladelphia|0.0|0.0|1.0|0.0|Woman Who Got Married in Blizzard Votes With Newborn Girl https://t.co/PLPAXbjbCO
AliciaBarnesTV|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
AliciaBarnesTV|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
ruchdesh|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
BubashLance|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
JeromeChallamel|SkyNews|0.0|0.0|1.0|0.0|Also Live #ElectionResults via @SkyNews https://t.co/M6rpVJ94Z8 #Election2016 #ElectionDay #ElectionNight #HillaryClinton #DonaldTrump
JeromeChallamel|election|0.0|0.0|1.0|0.0|Also Live #ElectionResults via @SkyNews https://t.co/M6rpVJ94Z8 #Election2016 #ElectionDay #ElectionNight #HillaryClinton #DonaldTrump
iJasonYu|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
iJasonYu|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
209twitch|MaxMeleganich|-0.1531|0.348|0.652|0.0|@MaxMeleganich @inshaIlah awkward https://t.co/4vRGCllGBU
209twitch|nytimes|-0.1531|0.348|0.652|0.0|@MaxMeleganich @inshaIlah awkward https://t.co/4vRGCllGBU
mrn9b|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
OmarMR709|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
OmarMR709|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
u2_lisa|tonygoldwyn|0.7772|0.0|0.702|0.298|@tonygoldwyn Tony Goldwyn!!! Are you ready to make history?! Never been so excited about an election! #ElectionNight https://t.co/9pX7vSCj25
u2_lisa|twitter|0.7772|0.0|0.702|0.298|@tonygoldwyn Tony Goldwyn!!! Are you ready to make history?! Never been so excited about an election! #ElectionNight https://t.co/9pX7vSCj25
ericathas|npr|0.0|0.0|1.0|0.0|The @npr live blog--&gt; https://t.co/IYdhOSnhEqState-by-state results--&gt; https://t.co/qx1CdIqJafContext--&gt; https://t.co/EatqgPk7XL
ericathas|t|0.0|0.0|1.0|0.0|The @npr live blog--&gt; https://t.co/IYdhOSnhEqState-by-state results--&gt; https://t.co/qx1CdIqJafContext--&gt; https://t.co/EatqgPk7XL
Karl_Huebner|tomjensen100|-0.34|0.146|0.854|0.0|RT @tomjensen100: This election has me stressed out. May be time for a Mazel Tov Cocktail.
ASUCRiverside|facebook|0.0|0.0|1.0|0.0|Fellow #Highlanders! Tonight there will be a live Election Coverage event in HUB 302! This is a historical... https://t.co/mBThJmwNih
JustinWelham|CharlieDayQuote|0.0|0.0|1.0|0.0|RT @CharlieDayQuote: After the election results tonight... https://t.co/cmPwW4Jded
JustinWelham|twitter|0.0|0.0|1.0|0.0|RT @CharlieDayQuote: After the election results tonight... https://t.co/cmPwW4Jded
worldnews_net|abcnews|0.0|0.0|1.0|0.0|How Donald Trump Is Spending Election Night https://t.co/zmNZ6HvF1w #abcnews #abc #news
annie773|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
BernThe270|twitter|0.0|0.0|1.0|0.0|ELECTION PROTECTION#API Asian Pacific IslanderAAJC's #VoterHotline for non-English speakers.800-API-VOTE https://t.co/wRJdCic8n3
TroyChildress1|vfmeadows17|0.5719|0.0|0.709|0.291|RT @vfmeadows17: Happy Election Day franz  #MAGA #TrumpTrain @OldRowOfficial https://t.co/65pMbrLUpe
TroyChildress1|twitter|0.5719|0.0|0.709|0.291|RT @vfmeadows17: Happy Election Day franz  #MAGA #TrumpTrain @OldRowOfficial https://t.co/65pMbrLUpe
malindalo|instagram|0.0|0.0|1.0|0.0|Election night apple galette! #homecooking #baking https://t.co/mdUtwPBIzb
SmallFriesBaby|tyleroakley|0.861|0.0|0.687|0.313|"RT @tyleroakley: better late than never!! if you've never voted before, make THIS election your first. it's so easy &amp; you won't regret it."
saintjada13|kelly_ohmann|-0.624|0.281|0.611|0.108|RT @kelly_ohmann: if I have to hear one more privileged ass white boy say this election doesn't matter I am going to LOSE IT
doctor_oddball|jimsciutto|0.0|0.0|1.0|0.0|"@jimsciutto @Stefan_Laurell @KristinFisher They should have taken a ""nutscape"" photo of earth for this election"
kanimozhi|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
GOPbattle2016|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
autobody65|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
lucy__hannah__|CallmeQueen_G|-0.3612|0.179|0.718|0.103|"RT @CallmeQueen_G: Plot twist: this whole election was a bad dream, and Bernie Sanders is actually president"
acpcsn|voxdotcom|0.0|0.0|1.0|0.0|"Pantsuit Nation, the giant, secret Hillary Facebook group, explained https://t.co/MK06IlwK3A via @voxdotcom"
acpcsn|vox|0.0|0.0|1.0|0.0|"Pantsuit Nation, the giant, secret Hillary Facebook group, explained https://t.co/MK06IlwK3A via @voxdotcom"
garryshown|mike_pence|0.3818|0.0|0.894|0.106|"RT @mike_pence: The outcome of this historic election rests in your hands. If you stand for a stronger America, cast your vote for #TrumpPe"
noropthony|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
CarlosHerrera|inti|0.0|0.0|1.0|0.0|RT @inti: President | Live Election Night Forecast | FiveThirtyEight https://t.co/8Lqe5XUdrA #ElectionDay
CarlosHerrera|projects|0.0|0.0|1.0|0.0|RT @inti: President | Live Election Night Forecast | FiveThirtyEight https://t.co/8Lqe5XUdrA #ElectionDay
bianca_mansour|marcieyounis|0.5859|0.0|0.703|0.297|RT @marcieyounis: the real winner of the presidential election. https://t.co/bBCIF6MGeF
bianca_mansour|twitter|0.5859|0.0|0.703|0.297|RT @marcieyounis: the real winner of the presidential election. https://t.co/bBCIF6MGeF
Mendoza11A|CJ_Squad11|0.0|0.0|1.0|0.0|RT @CJ_Squad11: Realist Thing About Today's Election. https://t.co/U2BgDu3H2I
Mendoza11A|twitter|0.0|0.0|1.0|0.0|RT @CJ_Squad11: Realist Thing About Today's Election. https://t.co/U2BgDu3H2I
dhcalalily28|DonaldJTrumpJr|0.3164|0.0|0.906|0.094|RT @DonaldJTrumpJr: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERSGET OUT AND VOTE! Find 5 others. This is our chance to take back Am
reblatt|kevindale|0.0|0.0|1.0|0.0|RT @kevindale: First live election show of the night about to start @cronkitenews https://t.co/YwMIVqqmAA
reblatt|twitter|0.0|0.0|1.0|0.0|RT @kevindale: First live election show of the night about to start @cronkitenews https://t.co/YwMIVqqmAA
halomoma|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
worldnews_net|latimes|0.0|0.0|1.0|0.0|Former President George W. Bush didn't vote for Donald Trump https://t.co/1CVbfh9MRJ #LosAngelesTimes #latimes #news
Red4Jacob|FailGOP|0.6369|0.0|0.781|0.219|RT @FailGOP: Might be one of the best things I have heard this entire election cycle. https://t.co/dcmTKGbUGM
Red4Jacob|twitter|0.6369|0.0|0.781|0.219|RT @FailGOP: Might be one of the best things I have heard this entire election cycle. https://t.co/dcmTKGbUGM
tcolkos98|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
taliadelrey|THOTJAI|0.5719|0.0|0.821|0.179|RT @THOTJAI: if donald trump wins the election I will paypal 100 dollars to everyone that retweets this #ElectionDay
goodforsumthin|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: Ohio, it's Election Day! Polls are open from 6:30am-7:30pm. Confirm your polling place now and go vote for Hillary! htt"
Lawgotsoul|CNNPolitics|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
Lawgotsoul|twitter|0.0|0.0|1.0|0.0|RT @CNNPolitics: Stand by for #CNNElection projectionhttps://t.co/jOauYyVeuX#ElectionNight https://t.co/8Jx61W8ceh
DenniLeigh|LJSRileyJohnson|0.0|0.0|1.0|0.0|"RT @LJSRileyJohnson: Voter ID is not required in almost all voter situations in NE, except in rare case detailed here by @NebraskaReform: h"
Basilswiss|twitter|-0.6115|0.154|0.846|0.0|"She must think a lot of people really hate her, and she hasn't even been elected yet. Wonder what she will do after https://t.co/kl8YjEvA9p"
TheScream666|mtv|0.0|0.0|1.0|0.0|333333333433333: RT MTVNews: wyd tonight? come thru 6:50pm ET  https://t.co/6rfZkhyZqB https://t.co/zM4JZ2axAP
galaxietoots|caribeauchamp|0.4215|0.0|0.877|0.123|RT @caribeauchamp: Off to Nancy Olson's to #nastywomenunite  After years of getting each other thru debates and election nights hoping for
thewickedlilith|CurveMe|0.6633|0.0|0.772|0.228|RT @CurveMe: IF TRUMP WINS THE ELECTION   IM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICAGOODMORNINGSAN DIEGO
donstanley72|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
donstanley72|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
TheBlindDonkey|PasadenaNow|0.8122|0.0|0.654|0.346|Thanks to @PasadenaNow for naming us one of the best places to drink after voting!https://t.co/LKUHaT9UVq https://t.co/pNDLhkR07a
TheBlindDonkey|pasadenanow|0.8122|0.0|0.654|0.346|Thanks to @PasadenaNow for naming us one of the best places to drink after voting!https://t.co/LKUHaT9UVq https://t.co/pNDLhkR07a
TheSaintKopite|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
TheSaintKopite|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
the_herald|TheBlogDH|0.0|0.0|1.0|0.0|RT @TheBlogDH: Big day for election coverage! We will be live blogging and on Facebook/Twitter throughout the night as our next president i
yaydal|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
accumulationwp|fivethirtyeight|0.2023|0.0|0.899|0.101|How important is Florida? (Polls in the eastern part of the stateclose in a few minutes.) If https://t.co/iH1uMyoVxl
summerleyphoto|DannyAustin_9|0.0|0.0|1.0|0.0|"RT @DannyAustin_9: Folks already getting seats for election results in Times Square, according to one dude ... Six hours before polls close"
Gfabgab|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Gfabgab|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
joeyalison|twitter|-0.8779|0.359|0.641|0.0|"Me just now: Oh, fuck, what the fuck is this election map, oh jesus...wait, this is a goddamn cell phone ad. https://t.co/hy3EPXLCyw"
_CHRIS__Cross|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
DaisyHavoc|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
63_DTiger|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
63_DTiger|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
Izengabe_|RRHElections|0.0|0.0|1.0|0.0|"RT @RRHElections: Our liveblog is, err, live! Starting in Kentucky, working our way up to Indiana. https://t.co/sv9zuGjp8Q"
Izengabe_|rrhelections|0.0|0.0|1.0|0.0|"RT @RRHElections: Our liveblog is, err, live! Starting in Kentucky, working our way up to Indiana. https://t.co/sv9zuGjp8Q"
itsmemaggieno7|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
itsmemaggieno7|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
daRude83|SenBernie|-0.4086|0.242|0.64|0.118|Lets not forget the biggest loser of the election: @SenBernie #electionday
BrookLassie|twitter|-0.7995|0.353|0.479|0.168|TOTALLY illegal.  hillary cheated in debate why wouldn't she steal an election? The woman had NO interest at her ra https://t.co/41jRUujXDG
nicknow|instagram|0.6369|0.0|0.704|0.296|Political junkie...I love election night and now I don't have to https://t.co/kSYtSil6m2
UnkelFred|larochecbc|-0.6124|0.295|0.591|0.114|RT @larochecbc: As a Cdn watching US election. Feels like that slow drive past horrendous crash scene.
Lucashigdon24|Things4WhitePpl|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
Lucashigdon24|twitter|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
12wollmana|michaelianblack|-0.0516|0.132|0.746|0.123|RT @michaelianblack: Quick reminder that Paul Ryan and nearly the entire Republican leadership disgraced themselves at every opportunity th
athirahchan|thephilacitizen|-0.4019|0.119|0.881|0.0|"RT @thephilacitizen: We've teamed with @votecastr for live voting results all day. Now, Clinton leading in the first battleground state: ht"
dman11235|dman11235|-0.802|0.313|0.687|0.0|@dman11235 The problem is that it came out a week ago that his competition literally broke election laws.  He'll lose by 2 points.
doparrish51|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
doparrish51|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
morgan__joy|TheQueenTee_|-0.4767|0.256|0.744|0.0|RT @TheQueenTee_: our nation is crying over this election https://t.co/bzE1ficzqI
morgan__joy|twitter|-0.4767|0.256|0.744|0.0|RT @TheQueenTee_: our nation is crying over this election https://t.co/bzE1ficzqI
amcomis|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
amcomis||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
bamamom2x|yankeebrit77|0.0|0.0|1.0|0.0|@yankeebrit77 @redostoneage Soros election rigging software and machines!
dmillerwats|CNN|0.3182|0.0|0.881|0.119|RT @CNN: Warren Buffett has kept his promise to drive voters to the polls on #ElectionDay https://t.co/qJZl9WZhRH https://t.co/7vhuoGlqdQ
dmillerwats|money|0.3182|0.0|0.881|0.119|RT @CNN: Warren Buffett has kept his promise to drive voters to the polls on #ElectionDay https://t.co/qJZl9WZhRH https://t.co/7vhuoGlqdQ
Time_New_Marcus|Battlefieldtrip|0.3612|0.0|0.865|0.135|RT @Battlefieldtrip: I've got my 2017 style on lock - are YOU ready for the post-election wasteland? https://t.co/sC0Sf5Gw7V
Time_New_Marcus|twitter|0.3612|0.0|0.865|0.135|RT @Battlefieldtrip: I've got my 2017 style on lock - are YOU ready for the post-election wasteland? https://t.co/sC0Sf5Gw7V
Paul55770744|linkis|0.9114|0.0|0.527|0.473|SEE IT! Madonna withdraws oral sex promise to Hillary voters https://t.co/nFe5tnhgGn. HA HA HA!! Have to watch video
payneywayney7|CNNPolitics|0.0|0.0|1.0|0.0|RT @CNNPolitics: The first polls are closing at 7 p.m. ET. Get the latest results here https://t.co/jOauYyVeuX https://t.co/inPimatat2
payneywayney7|cnn|0.0|0.0|1.0|0.0|RT @CNNPolitics: The first polls are closing at 7 p.m. ET. Get the latest results here https://t.co/jOauYyVeuX https://t.co/inPimatat2
mel_huang|politico's|0.1779|0.145|0.633|0.222|"Ok, clearly @politico's election maps are not working right and they do not have updated data. Disappointing."
jesdaleo|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
MattPosorske|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
SirDickOfHearts|tinkersong|-0.4588|0.15|0.85|0.0|@tinkersong I think both should be banned from covering any election once the polls open and until they close.
fangpusskins|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
fangpusskins|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
TheAtomicRaygun|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
t045tbr0t|Suxting|0.3182|0.0|0.685|0.315|RT @Suxting: I've got a huge election.
krazyjake313|mike_pence|0.0|0.0|1.0|0.0|"RT @mike_pence: This Election Day, America is standing at the crossroads of history. RT this if you're voting for @realDonaldTrump. Togethe"
_Proud_American|bunkerwsmith|0.5574|0.063|0.704|0.233|"RT @bunkerwsmith: To people feeling anxiety about the election: Focus on things you can control, like VOTING. Keep your chin up. Stay calm."
highkeyme_|twitter|0.0|0.0|1.0|0.0|Very appropriate tweet for this election!  https://t.co/rTrWeUFVVq
abern918|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
TheSteeldawn|Khaixur|-0.743|0.259|0.741|0.0|"@Khaixur If it's proven that clinton rigged states with voter fraud and election rigs, then trump ends up being right."
TweetieDede|twitter|0.6887|0.0|0.77|0.23|Stay tuned for a key Tweetie Dede election night alert ... Not really just laughing at the pundits early time fille https://t.co/xe6xuQYtCU
quiddlet|twitter|0.0|0.0|1.0|0.0|Took until election day but the metaphor is complete. https://t.co/K7QUYSHYQ4
KristaGuida|instagram|0.4939|0.0|0.824|0.176|"I know, I know, there's an election and SUCH exciting talk and speculation for HOURS about who https://t.co/d3rVHjWaBf"
worldnews_net|latimes|0.0|0.0|1.0|0.0|How this election has revealed workplace sexism is still an issue https://t.co/jH1iqRWNbJ #LosAngelesTimes #latimes #news
MRODDDY|MelisaFranzen|0.0|0.0|1.0|0.0|Hitting the doors one last time for @MelisaFranzen on election night! THIS is how we make a change. THIS is how we https://t.co/wEPms2ysk8
MRODDDY|twitter|0.0|0.0|1.0|0.0|Hitting the doors one last time for @MelisaFranzen on election night! THIS is how we make a change. THIS is how we https://t.co/wEPms2ysk8
Zachendowed|Derek74399105|-0.6253|0.212|0.788|0.0|"RT @Derek74399105: The American election is very dull and not rossy like Nigeria election , nobody snatch ballot box, agbero didn't break"
notime2write|Isaacsvillegas|0.5719|0.0|0.773|0.227|RT @Isaacsvillegas: Leftover Halloween candy. Vital for Election Day. I recommend the funsize snickers bars. Healthiest because peanuts. #s
ScottMitch77|EW|0.4019|0.0|0.828|0.172|"https://t.co/xxkcSKlEHu: ""Laura Benanti appearing on Stephen Colbert's election night special on Showtime"" @EW https://t.co/vUhYSge4Sm"
ScottMitch77|ew|0.4019|0.0|0.828|0.172|"https://t.co/xxkcSKlEHu: ""Laura Benanti appearing on Stephen Colbert's election night special on Showtime"" @EW https://t.co/vUhYSge4Sm"
throbbjon|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
blujaydavid|PerezHilton|0.0|0.0|1.0|0.0|RT @PerezHilton: #HillaryClinton does the #MannequinChallenge for #ElectionDay! https://t.co/EBHYc5eVrt https://t.co/i5Dz7zPnDo
blujaydavid|perezhilton|0.0|0.0|1.0|0.0|RT @PerezHilton: #HillaryClinton does the #MannequinChallenge for #ElectionDay! https://t.co/EBHYc5eVrt https://t.co/i5Dz7zPnDo
pedrobroa|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/GoYnDeEvaH
pedrobroa|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/GoYnDeEvaH
randomsweede|LeahR77|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
randomsweede|breitbart|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
SHAEkeIt_Baby|yupDESme_|0.0|0.0|1.0|0.0|RT @yupDESme_: someone explain to me why high schoolers get out of school for Election Day but college students..that can actually vote..st
L0Lbasic|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
justjaney_|korndiddy|0.2561|0.0|0.904|0.096|RT @korndiddy: So... you're telling me I'm expected to do actual work today? ...And not just anxiously refresh election news?
janakatharine8|hollywoodreporter|0.6369|0.0|0.543|0.457|Hollywood's best #Election2016 tweets https://t.co/l5IkIvyExH https://t.co/KJDYPckY8g
reisegrrl1|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
UrbanismAvenger|ajplus|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
UrbanismAvenger|twitter|-0.5574|0.195|0.805|0.0|RT @ajplus: Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/uHRaxDceau
BrandonLRichard|ABC|0.0|0.0|1.0|0.0|RT @ABC: ELECTION NIGHT: Who will be our next president? Coverage starting at 7PM ET on @ABCNetwork and across @ABC digital: https://t.co/V
BrandonLRichard|t|0.0|0.0|1.0|0.0|RT @ABC: ELECTION NIGHT: Who will be our next president? Coverage starting at 7PM ET on @ABCNetwork and across @ABC digital: https://t.co/V
emeraldfury|heraldleader|0.0|0.0|1.0|0.0|RT @heraldleader: Updating state House results: https://t.co/96mFP7TyEd https://t.co/sFQZSDXGvY
emeraldfury|kentucky|0.0|0.0|1.0|0.0|RT @heraldleader: Updating state House results: https://t.co/96mFP7TyEd https://t.co/sFQZSDXGvY
MrEdTrain|surfermom77|0.0|0.0|1.0|0.0|"RT @surfermom77: Twitter &amp; FB R begin inundated wt reports of Elec.fraud, voting irregularities &amp; discrimination against Trump Votershttps"
LonelyLizards|YouTube|0.0|0.0|1.0|0.0|election day: https://t.co/RPUx25gZPr via @YouTube
LonelyLizards|youtube|0.0|0.0|1.0|0.0|election day: https://t.co/RPUx25gZPr via @YouTube
Mr3lsewhere|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
Mr3lsewhere|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
tony_ganzer|NickCastele|0.0|0.0|1.0|0.0|RT @NickCastele: Director of @cuyahogaboe says rumored self-appointed Trump election observers didn't show up at polling places here.
caligramma|EricBoehlert|0.5574|0.0|0.783|0.217|RT @EricBoehlert: we should rename Election Day to Laugh At James O'Keefe Day https://t.co/q7EPl32Zly
caligramma|twitter|0.5574|0.0|0.783|0.217|RT @EricBoehlert: we should rename Election Day to Laugh At James O'Keefe Day https://t.co/q7EPl32Zly
deejjaaj|piercespears|0.5719|0.0|0.829|0.171|RT @piercespears: Historians will look back at this video and say this is why Hillary won the election  https://t.co/aaAKHIKPyv
deejjaaj|twitter|0.5719|0.0|0.829|0.171|RT @piercespears: Historians will look back at this video and say this is why Hillary won the election  https://t.co/aaAKHIKPyv
ottdogbuns|Suxting|0.3182|0.0|0.685|0.315|RT @Suxting: I've got a huge election.
sarsoorra|G_Eazy|0.7644|0.0|0.752|0.248|"RT @G_Eazy: PLEASE GO OUT AND VOTE WHATEVER YOU DO, THIS COULD BE THE MOST IMPORTANT ELECTION OF OUR LIVES #imwithher #fuckdonaldtrump"
anthonyzupa|onsomeshit|-0.296|0.109|0.891|0.0|RT @onsomeshit: CNN just interrupted their election coverage to report on @lilyachty not knowing the words to Big Poppa
buckitman|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
BlastingNews|us|0.0|0.0|1.0|0.0|#election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR https://t.co/AfJAdNdbSU
efairhurst|vogue|0.0|0.0|1.0|0.0|Daniel Arnold Talks Politics With New York City Voters on Election Day https://t.co/IAmhCiu0OS
Avocadohomo|lntroset|0.8969|0.0|0.67|0.33|RT @lntroset: Today is Election Day so I thought I would share the loving someone lyrics with you guys bc this world needs more love and le
ddhorn4065|ananavarro|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
ddhorn4065|twitter|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
jakeroberts2015|YahooNews|-0.8689|0.353|0.647|0.0|RT @YahooNews: WATCH LIVE: GOP pollster @FrankLuntz says Its a vote between a liar and a lunatic &amp; people will choose the liar https://t
jakeroberts2015||-0.8689|0.353|0.647|0.0|RT @YahooNews: WATCH LIVE: GOP pollster @FrankLuntz says Its a vote between a liar and a lunatic &amp; people will choose the liar https://t
JeffroJoiner|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
JeffroJoiner|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
rabuliz|DonaldJTrumpJr|0.8439|0.062|0.62|0.318|RT @DonaldJTrumpJr: No excuse not to vote. It is your duty to do everything you can to help save America. We can win this thing! #MAGA #Ele
biasbreakdown|NickTimiraos|-0.296|0.109|0.891|0.0|"RT @NickTimiraos: When the AP called the election2012: 11:38 pm, Tuesday2008: 11 pm, Tuesday2004: 11:19 am, Wednesday2000: No call1996"
kiaraxcook|gaileyfrey|0.3412|0.0|0.909|0.091|RT @gaileyfrey: Can you guys imagine if you were a little duckling right now If you didn't have to worry about the election &amp; could just
tabfishsg|JenJFielding|-0.6808|0.219|0.781|0.0|"RT @JenJFielding: Everyone's freaking out about the election, and I'm over freaking out about the new graphic design updates coming to #Tab"
margare79163346|LeeCamp|0.0|0.0|1.0|0.0|RT @LeeCamp: How do YOU feel about this #election?? #ElectionDay #Elections2016
jessjeffries1|Maddynx|0.0|0.0|1.0|0.0|RT @Maddynx: Twitter on Election Dayhttps://t.co/04p0nkjyiw
faobobindc|Kevin_Harron|0.0|0.0|1.0|0.0|RT @Kevin_Harron: Does @MSNBC put steve kornacki in a utility closet along with his magic election board until the next election after toni
TonyRocha__|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
TonyRocha__|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
GonnaRememberMe|hiimariela|0.6299|0.061|0.697|0.242|RT @hiimariela: so like after election is done who's down to take shots i need to calm all my nerves
THE_REAL_DESPO|Jerradjrod25|0.5598|0.0|0.795|0.205|RT @Jerradjrod25: @THE_REAL_DESPO trooooof fam so true all talking bout puppet election got me https://t.co/3SBt09s6cp
THE_REAL_DESPO|twitter|0.5598|0.0|0.795|0.205|RT @Jerradjrod25: @THE_REAL_DESPO trooooof fam so true all talking bout puppet election got me https://t.co/3SBt09s6cp
bitchywaiter|facebook|0.0|0.0|1.0|0.0|"Now, as we begin to watch election returns, a moment of silence for the livers that so many of us will lose... https://t.co/j2vWyhFNVK"
ElizabethClyde|MattBellassai|-0.25|0.264|0.566|0.17|RT @MattBellassai: my top Election Day worries: https://t.co/Qs3dIGh8uT
ElizabethClyde|twitter|-0.25|0.264|0.566|0.17|RT @MattBellassai: my top Election Day worries: https://t.co/Qs3dIGh8uT
DFSRotoMonsters|mikeeaves|0.0|0.0|1.0|0.0|"RT @mikeeaves: While Election2016 #ExitPolls Expected At 5PM EST, Here Is A Poll Closing Map To Follow The Actual Election Returns: https:/"
DFSRotoMonsters||0.0|0.0|1.0|0.0|"RT @mikeeaves: While Election2016 #ExitPolls Expected At 5PM EST, Here Is A Poll Closing Map To Follow The Actual Election Returns: https:/"
Love_Chihuahua|astroterf|0.0|0.0|1.0|0.0|RT @astroterf: Every election it's the SOS. WTF?! https://t.co/z38UNyzYJ4
Love_Chihuahua|twitter|0.0|0.0|1.0|0.0|RT @astroterf: Every election it's the SOS. WTF?! https://t.co/z38UNyzYJ4
pizdapalace|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
beckybazjones||0.3818|0.094|0.667|0.239|Alright everyone:  Solution to the anxiety of election results... Tuesday $5.00 movies @ Marcus Theatre. #letsgo
NBCNewYork|nbcnewyork|0.6124|0.0|0.583|0.417|These kindergartners just won the mannequin challenge https://t.co/d4RXMUnNXs https://t.co/RljwEfQ7Yd
mauisrf7|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
mauisrf7|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
jmsexton_|motherjones|0.0|0.0|1.0|0.0|It's Election Day and Fox News Just Had a Total Meltdown https://t.co/kzEvKlubLY  MoJo #ImWithHer #UniteBlue https://t.co/BN3ONjlNvL
krystalvivian|instagram|0.0|0.0|1.0|0.0|Election Night Pizza is the real MVP https://t.co/KM2i1id74T https://t.co/UZx1HrCy70
shernandez227|themoneygame|0.5719|0.0|0.821|0.179|RT @themoneygame: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/RTr54mdgR3 https://t.co/y
shernandez227|businessinsider|0.5719|0.0|0.821|0.179|RT @themoneygame: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/RTr54mdgR3 https://t.co/y
bbs_firstfed|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
GeorgiaDaskalos|DRUDGE_REPORT|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
GeorgiaDaskalos|businessinsider|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
psuba98|EveryonesLocal|-0.4019|0.13|0.81|0.061|RT @EveryonesLocal: Feeling masochistic? Come &amp; watch the  election results w us tonite on big screens - find out tonite if we need borde
rollecoarster|DanaiGurira|0.783|0.0|0.567|0.433|RT @DanaiGurira: Happy Election Day!Make sure your voice is heard!Vote!#ImWithHer.#TheFutureisFemale https://t.co/s6XK0ZYDzt
rollecoarster|twitter|0.783|0.0|0.567|0.433|RT @DanaiGurira: Happy Election Day!Make sure your voice is heard!Vote!#ImWithHer.#TheFutureisFemale https://t.co/s6XK0ZYDzt
AlanmBeat|WDFx2EU8|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
AlanmBeat|conservativeeagles|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
CherifLoutfi|YouTube|0.0|0.0|1.0|0.0|For those who are interrested  Decision 2016: LIVE Election Night Coverage | NBC News https://t.co/YUyrqM5uU6 via @YouTube
CherifLoutfi|youtube|0.0|0.0|1.0|0.0|For those who are interrested  Decision 2016: LIVE Election Night Coverage | NBC News https://t.co/YUyrqM5uU6 via @YouTube
CallHerAshley|paulafaris|0.4019|0.0|0.863|0.137|"RT @paulafaris: Here. We. Go. Gearing up for our @ABCNews election special, anchored by @GStephanopoulos and @MarthaRaddatz. https://t.co/J"
CallHerAshley|twitter|0.4019|0.0|0.863|0.137|"RT @paulafaris: Here. We. Go. Gearing up for our @ABCNews election special, anchored by @GStephanopoulos and @MarthaRaddatz. https://t.co/J"
Koxinga8|breitbart|0.0516|0.145|0.699|0.156|Nate Silver: Polling Error Could Be 'Higher Than Usual' Thanks to Late-Breaking Undecideds - Breitbart https://t.co/1eKn4TIHfH
cellydoumerc|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
siannelson1|sbrownson10|0.6369|0.0|0.826|0.174|RT @sbrownson10: Love how America is waiting for the presidential election and we're waiting to watch celebrities eat kangaroo bollocks aga
blueefoxxx|mikethenice1|0.0|0.0|1.0|0.0|"RT @mikethenice1: As The Election Comes To A Close, Turnout At Trump Rallies Is Massive https://t.co/wfwytJir8F"
blueefoxxx|westernjournalism|0.0|0.0|1.0|0.0|"RT @mikethenice1: As The Election Comes To A Close, Turnout At Trump Rallies Is Massive https://t.co/wfwytJir8F"
emuhlyyx3|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
PCNHCarey|twitter|0.0|0.0|1.0|0.0|Election pizza has arrived! #BayVotes https://t.co/u1Ov4QfEbm
The_Yodacat|KedgeOnline|0.0|0.0|1.0|0.0|"@KedgeOnline Turns out, the election was inside of us all along."
carlyburdett|SidneyCrosbyEgo|0.765|0.0|0.752|0.248|RT @SidneyCrosbyEgo: The best part about election day is that we get to watch McDavid and Crosby play before the world ends.
remzelk1|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
iShygga|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
iShygga|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
worldnews_net|latimes|0.0|0.0|1.0|0.0|"In Little Saigon, a possible generational divide at the polls https://t.co/sVw8Um6STb #LosAngelesTimes #latimes #news"
ghawtho1|OPB|-0.3818|0.148|0.852|0.0|"RT @OPB: At Susan B. Anthony's Grave, visiting hours extended for election day crowds  https://t.co/KWJS1XealL https://t.co/YItRaU3xO1"
ghawtho1|opb|-0.3818|0.148|0.852|0.0|"RT @OPB: At Susan B. Anthony's Grave, visiting hours extended for election day crowds  https://t.co/KWJS1XealL https://t.co/YItRaU3xO1"
265961fc22994f5|politico|0.0|0.0|1.0|0.0|"RT @politico: #BREAKING: Results of the U.S. elections are beginning to flow in, starting with returns from Indiana and Kentucky https://t."
265961fc22994f5||0.0|0.0|1.0|0.0|"RT @politico: #BREAKING: Results of the U.S. elections are beginning to flow in, starting with returns from Indiana and Kentucky https://t."
BarbaraB777|terrysumpter|-0.6166|0.335|0.665|0.0|RT @terrysumpter: OBAMA HAS FAILED AMERICA https://t.co/Vy2jzx6BRj via @BreitbartNews
BarbaraB777|breitbart|-0.6166|0.335|0.665|0.0|RT @terrysumpter: OBAMA HAS FAILED AMERICA https://t.co/Vy2jzx6BRj via @BreitbartNews
ss396camaro|0hour|0.0|0.0|1.0|0.0|RT @0hour: https://t.co/2S72Q1xk2DIndiana70% as of nowits happening!
ss396camaro|t|0.0|0.0|1.0|0.0|RT @0hour: https://t.co/2S72Q1xk2DIndiana70% as of nowits happening!
jamieraegomes|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
jamieraegomes|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
Danny_Bermudez|BuzzFeed|-0.6249|0.227|0.773|0.0|This is the worst content ever for election night. Get a new team @BuzzFeed @BuzzFeedNews #ElectionNight
HermanMcflurman|nytopinion|-0.34|0.111|0.841|0.049|RT @nytopinion: This election WAS rigged  by state governments that did all they could to prevent nonwhite Americans from voting. https://
HermanMcflurman||-0.34|0.111|0.841|0.049|RT @nytopinion: This election WAS rigged  by state governments that did all they could to prevent nonwhite Americans from voting. https://
Jesmeshd94|WORLDSTAR|0.5859|0.0|0.678|0.322|RT @WORLDSTAR: Who will win the 2016 presidential election? 
Tigresauce|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
Tigresauce|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
sri9011|smarket|-0.2732|0.091|0.909|0.0|RT @smarket: Modi should now follow this up by slashing Income Tax to 10% for income upto 10 lakhs...next election in bag
WSJ|WSJPolitics|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
WSJ|wsj|-0.3818|0.133|0.867|0.0|"RT @WSJPolitics: People line up to visit Susan B. Anthony's grave in Rochester, N.Y. on #ElectionDay https://t.co/svBB8C8bLY  https://t.co"
karenfeagins|teamvincek|0.5994|0.0|0.811|0.189|RT @teamvincek: Join @WJCTJax &amp; @NPR for live coverage of #ElectionNight. Tune in on 89.9 FM at 7 p.m. for our election special  https://t.
karenfeagins||0.5994|0.0|0.811|0.189|RT @teamvincek: Join @WJCTJax &amp; @NPR for live coverage of #ElectionNight. Tune in on 89.9 FM at 7 p.m. for our election special  https://t.
ProblematicRec|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
pacificgio|SebGorka|0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
pacificgio||0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
ph3ezus|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
analyticalps|DeplorableDJT|0.0|0.0|1.0|0.0|"@DeplorableDJT @NRO @marcorubio can we focus on this election, FIRST!"
jeanne_tall|Hardline_Stance|-0.9124|0.493|0.507|0.0|"RT @Hardline_Stance: massive VOTER FRAUD in #FTL #FL; Election workers caught faking 1,000's of stolen absentee ballotshttps://t.co/0ajn3"
SpinnakerPix|fivethirtyeight|0.0|0.0|1.0|0.0|I'm putting my money on @fivethirtyeight this #election
drkateyun|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
newspalmique|foxnews|0.0|0.0|1.0|0.0|#LatestNews LIVE COVERAGE Watch Fox News Channel Election Day 2016 coverage https://t.co/DAXeTGmTC4 by @foxnews
newspalmique|video|0.0|0.0|1.0|0.0|#LatestNews LIVE COVERAGE Watch Fox News Channel Election Day 2016 coverage https://t.co/DAXeTGmTC4 by @foxnews
actindia|DipDhingani|0.9091|0.0|0.55|0.45|"RT @DipDhingani: #Trump might win the election, but #Modi won the hearts. Haha. #blackmoney #FightAgainstCorruption #OnThisDay #CurrencyB"
Legochanful|GameTheoryRejct|-0.2323|0.193|0.652|0.155|RT @GameTheoryRejct: Meta Theory: Donald Trump will win the election WITH THE POWER OF THE CHAOS EMERALDS?! https://t.co/44jaJJ7Joq
Legochanful|twitter|-0.2323|0.193|0.652|0.155|RT @GameTheoryRejct: Meta Theory: Donald Trump will win the election WITH THE POWER OF THE CHAOS EMERALDS?! https://t.co/44jaJJ7Joq
jackodonnell96|JonErlichman|0.0|0.0|1.0|0.0|RT @JonErlichman: Things that didn't exist election night in 2008:UberiPadInstagramSnapchatWhatsAppPinterestPeriscopeOculusSlack
TonyBeavers1|LeahR77|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
TonyBeavers1|breitbart|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
AzadCandace|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
Hbkjoey2275|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
aineeyusry|AdaApaDgnCikTeh|0.7184|0.047|0.738|0.215|"RT @AdaApaDgnCikTeh: As much as CikTeh would love to joke about the American Election, I also have to take a hard look in the mirror to adm"
oldschoolvet74|viralnewsx|0.6523|0.1|0.651|0.249|"RT @viralnewsx: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://t.c"
oldschoolvet74||0.6523|0.1|0.651|0.249|"RT @viralnewsx: ELECTION DAY POLL: AFTER ALL THE MEDIA MANIPULATION AGAINST TRUMP, DO YOU BELIEVE HE STILL HAS A CHANCE TO WIN? https://t.c"
WinKox|CNN's|0.0|0.0|1.0|0.0|Watching @CNN's Election Night in America. #ElectionDay
sarahjaneb0rean|VP|0.0|0.0|1.0|0.0|RT @VP: Today is Election Day in America. Its time to get out and vote. https://t.co/a0MJUF4QIy
sarahjaneb0rean|twitter|0.0|0.0|1.0|0.0|RT @VP: Today is Election Day in America. Its time to get out and vote. https://t.co/a0MJUF4QIy
AidCourtney|SusanCalman|0.3612|0.0|0.848|0.152|RT @SusanCalman: Now for the election. I'm staying up all night.  I have provisions. I'm ready.
alexisbahl1603|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
DonkeyPunch145|twitter|-0.2732|0.231|0.769|0.0|Even ESPN is nervous about this election. https://t.co/XMZiJ4QX1S
GAFan8|JaimeeLiegh|-0.2732|0.123|0.877|0.0|RT @JaimeeLiegh: I don't even live in America and yet the election is making me nervous #ElectionNight
suz_stone|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
johnnyfire817|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
johnnyfire817|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
mannicmo2001|RT_America|-0.4019|0.153|0.847|0.0|"RT @RT_America: BREAKING: Polling station on lockdown after shooting leaves 2 injured in Azuza, CA https://t.co/G0cuZ0bfH0 https://t.co/ffi"
mannicmo2001|rt|-0.4019|0.153|0.847|0.0|"RT @RT_America: BREAKING: Polling station on lockdown after shooting leaves 2 injured in Azuza, CA https://t.co/G0cuZ0bfH0 https://t.co/ffi"
dcutler1958|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
dcutler1958|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
LifeOfNadom|boostmobile|0.4404|0.0|0.873|0.127|RT @boostmobile: 3.5 hr early voting wait in Los Angeles. Everyone deserves easy access to the polls. Sign below to #BoostYourVoicehttps:
bethanycarol1|ananavarro|0.9455|0.0|0.463|0.537|Thank you @ananavarro for your fierce passion- I have so enjoyed and admired your strong voice in this election!  https://t.co/npLHtAep4g
bethanycarol1|twitter|0.9455|0.0|0.463|0.537|Thank you @ananavarro for your fierce passion- I have so enjoyed and admired your strong voice in this election!  https://t.co/npLHtAep4g
gdsmack267|ESPNStatsInfo|0.34|0.0|0.906|0.094|RT @ESPNStatsInfo: Connor McDavid &amp; Sidney Crosby meet for 1st timeMario Lemieux &amp; Wayne Gretzky played vs each other for 1st time on Ele
gothdogs|twitter|0.4939|0.0|0.814|0.186|In honor of election night.....ask the gays what they think and what they do https://t.co/EHPg5sMj37
graywolf|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
PatriciaWilhoit|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
bedwcr|ladygaga|0.0|0.0|1.0|0.0|@ladygaga VOTE TRUMP. ONLY REAL PRESIDENT RUNNING THIS ELECTION.
Alex8awa|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
iceman120|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
jessicaseaman|alyrose|0.0|0.0|1.0|0.0|In the newsroom we have pizza for election night along with some cheese  dip   @alyrose https://t.co/Rq25rRo7zU
jessicaseaman|twitter|0.0|0.0|1.0|0.0|In the newsroom we have pizza for election night along with some cheese  dip   @alyrose https://t.co/Rq25rRo7zU
philmonaco67|WDFx2EU8|-0.1531|0.121|0.781|0.098|"RT @WDFx2EU8: The  election in a nutshell. On the left, Lady Gaga dancing like a dipshit at Clinton concert. On right, Mike Pence talking a"
Kilkenny_yyc|instagram|0.4574|0.0|0.857|0.143|"Red white and blue, America we are here for you! Kilkenny is having an election party and its https://t.co/KVlgl6QQ9X"
Bammers05|TBNSport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
Bammers05|tbnsport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
seaexpattrader|reuters|-0.6249|0.24|0.76|0.0|"First U.S. polls close as voters pick between Clinton, Trump after brutal campaign https://t.co/QW5L4qtijD"
bylaurenfitz|CPSuccessCHI|0.0|0.0|1.0|0.0|RT @CPSuccessCHI: .Brown: Student judges hold their own on Election Day #cpsuccess via @markbrowncst https://t.co/vhEiGn9725
bylaurenfitz|bit|0.0|0.0|1.0|0.0|RT @CPSuccessCHI: .Brown: Student judges hold their own on Election Day #cpsuccess via @markbrowncst https://t.co/vhEiGn9725
hoyawolf|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
hoyawolf|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
lisastokke|JamilSmith|-0.6486|0.249|0.751|0.0|"RT @JamilSmith: If it's Election Day, there are reports of voting disruptions. Machines malfunctioning, and people intimidating. https://t."
lisastokke||-0.6486|0.249|0.751|0.0|"RT @JamilSmith: If it's Election Day, there are reports of voting disruptions. Machines malfunctioning, and people intimidating. https://t."
Saeya8|immigrant4trump|0.7506|0.0|0.766|0.234|"RT @immigrant4trump: If you make this go viral, Trump will win. It's about 2 minutes that makes the choice in this election crystal clear h"
globalissuesweb|twib|0.0|0.0|1.0|0.0|America heads to the polls in 2016 elections  as it happened https://t.co/OysLeKsgiF https://t.co/iXgK8Cf0jQ
kungfujustice|MichaelHill51|0.1027|0.092|0.798|0.109|RT @MichaelHill51: The meaning of this election is clear: demographic warfare and the displacement of whites as a political force. This is
bobhardt|NY1|0.1779|0.122|0.718|0.16|An all-New York presidential election. No better place to watch all night long than @NY1
spnsammy|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
ricardowec|theverge|0.0|0.0|1.0|0.0|10 provocative political novels to read after the election https://t.co/VSaL5HGNaT #VergeNews
lhuffman34|vfmeadows17|0.5719|0.0|0.709|0.291|RT @vfmeadows17: Happy Election Day franz  #MAGA #TrumpTrain @OldRowOfficial https://t.co/65pMbrLUpe
lhuffman34|twitter|0.5719|0.0|0.709|0.291|RT @vfmeadows17: Happy Election Day franz  #MAGA #TrumpTrain @OldRowOfficial https://t.co/65pMbrLUpe
CityAndStateNY|JCColtin|0.0|0.0|1.0|0.0|"RT @JCColtin: Here at Javits for the Clinton election night event w/ @CityAndStateNY... and wifi is already slow! Gonna be a long, (hopeful"
notabasic_becca|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
wsjulian|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
wsjulian||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
josesolonh|ParisHilton|0.6094|0.0|0.801|0.199|RT @ParisHilton: This is one of the most important election's of our lifetime! Every vote makes a difference! Everyone please get out and #
lukescumstagram|1dsaints|0.6645|0.089|0.566|0.346|RT @1dsaints: please don't waste a vote. be smart about this election. this is not a joke https://t.co/m3hWDk3gEM
lukescumstagram|twitter|0.6645|0.089|0.566|0.346|RT @1dsaints: please don't waste a vote. be smart about this election. this is not a joke https://t.co/m3hWDk3gEM
bebebebender|Jonbuckhouse|0.6239|0.0|0.843|0.157|RT @Jonbuckhouse: The Polls are starting to close all over the US! Who do you think will win the election?  #ElectionNight #electionday #iV
9NewsMelb|9NewsAUS|0.0|0.0|1.0|0.0|"RT @9NewsAUS: .@LauraTurner_9 with Gary Langer, ABC News America Pollster, discussing how data is analysed. #ElectionDay #9News  https://t."
9NewsMelb||0.0|0.0|1.0|0.0|"RT @9NewsAUS: .@LauraTurner_9 with Gary Langer, ABC News America Pollster, discussing how data is analysed. #ElectionDay #9News  https://t."
rmcardz|0hour|0.0|0.0|1.0|0.0|RT @0hour: https://t.co/2S72Q1xk2DIndiana70% as of nowits happening!
rmcardz|t|0.0|0.0|1.0|0.0|RT @0hour: https://t.co/2S72Q1xk2DIndiana70% as of nowits happening!
allkbell|KathleenLights1|0.4199|0.141|0.573|0.286|RT @KathleenLights1: Hope everyone voted today! This election has traumatized me.... I pray for America.
mariajoseCANEL|nancybocskor|0.0|0.0|1.0|0.0|RT @nancybocskor: How I spent Election Day  550 people. 45 countries. https://t.co/28SsqeOZBs
mariajoseCANEL|twitter|0.0|0.0|1.0|0.0|RT @nancybocskor: How I spent Election Day  550 people. 45 countries. https://t.co/28SsqeOZBs
sylviagarner_|ItsWilliamD|0.0|0.0|1.0|0.0|"RT @ItsWilliamD: When autocorrect hits you with ""holy shot"".#lol #funny #harambe #ballislife #kenbone #memes #dankmemes #dank #tweet #jesu"
ohthatgizzmo|Impolitics|0.3182|0.0|0.913|0.087|"RT @Impolitics: This will always be remembered as the presidential election in which the KKK, the KGB and the FBI all supported the same ca"
smolkjd|NathanZed|-0.25|0.215|0.601|0.184|RT @NathanZed: I remember back when this election was all fun and games like when we accused a candidate of being a serial murderer can we
kfitz134|UNC_Humor|0.4404|0.0|0.791|0.209|"@UNC_Humor thanks to this election, our bell has never been more divided. "
KEVDSP10|SebGorka|0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
KEVDSP10||0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
thecimeshop|RT_America|-0.4019|0.153|0.847|0.0|"RT @RT_America: BREAKING: Polling station on lockdown after shooting leaves 2 injured in Azuza, CA https://t.co/G0cuZ0bfH0 https://t.co/ffi"
thecimeshop|rt|-0.4019|0.153|0.847|0.0|"RT @RT_America: BREAKING: Polling station on lockdown after shooting leaves 2 injured in Azuza, CA https://t.co/G0cuZ0bfH0 https://t.co/ffi"
SOgnenis|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
SOgnenis|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
LanzaJeremy|inzain98|0.4767|0.119|0.595|0.286|RT @inzain98: No matter who becomes President after this election I still love this country.
donna_grooms|TIME|-0.0258|0.073|0.927|0.0|RT @TIME: The overlooked history behind the movement to wear white on Election Day https://t.co/4aYW2SdOcG
donna_grooms|time|-0.0258|0.073|0.927|0.0|RT @TIME: The overlooked history behind the movement to wear white on Election Day https://t.co/4aYW2SdOcG
diasporaafro_|biggabossben|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
diasporaafro_|twitter|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
markagallolv|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: Drudge saying, ""Election will come down to evening voters.""  That means, ""Republicans with actual jobs."""
lezley_04|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
feministkraken|PatrioticSocks|0.0|0.0|1.0|0.0|"@PatrioticSocks @HullAmStuds @UniOfHull election night, @ualbany style! https://t.co/nY22fgqEw3"
feministkraken|twitter|0.0|0.0|1.0|0.0|"@PatrioticSocks @HullAmStuds @UniOfHull election night, @ualbany style! https://t.co/nY22fgqEw3"
JR777771|kindcutesteve|-0.5719|0.209|0.791|0.0|RT @kindcutesteve: MotherJones: This Election Is a Referendum on Hate (vote against it)#p2 #TNTweeters #USLatino #VoteBluehttps://t.co/Yj
TheMource|themource|0.2755|0.0|0.869|0.131|for more info https://t.co/6fXFivzEre Hillary Clinton -- Don't Mess W... https://t.co/nEp8eeyHqw #lol #cute #live https://t.co/EBi78lXDYa
SirLoinOBeef|FreddieCampion|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
SirLoinOBeef|twitter|0.6369|0.0|0.743|0.257|RT @FreddieCampion: Donald Trump makes good on his promise to have Election Day observers monitoring immigrants https://t.co/dRpDqhylzQ
TheReedsterr|everywordisgay|0.0|0.0|1.0|0.0|RT @everywordisgay: gay election
sammymoh|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
sammymoh|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
Jack_Eble_KDLT|KDLTNews|-0.5719|0.239|0.761|0.0|RT @KDLTNews: A fire incident at a Rapid City polling location will delay the results for #ElectionNight. #KDLTNews https://t.co/5jYgJxXXDs
Jack_Eble_KDLT|kdlt|-0.5719|0.239|0.761|0.0|RT @KDLTNews: A fire incident at a Rapid City polling location will delay the results for #ElectionNight. #KDLTNews https://t.co/5jYgJxXXDs
CurlyQEsq|conor64|-0.2411|0.073|0.927|0.0|RT @conor64: If you're still not sure whether you'll vote and you're waiting for a sign this is it: Go vote. This isn't the election to sit
ItsMattJordan|Glenn__Kenny|0.0|0.0|1.0|0.0|"RT @Glenn__Kenny: Remembering Election Day '80, when my Repub girlfriend took me to ""Sauve qui peut,"" a porn movie, &amp; ""Vampyr"" at Anthology"
Danieljackson94|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
Danieljackson94|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
AndyDavidJones|adubs_1|0.6369|0.0|0.811|0.189|"#Election2016 This just in... @adubs_1 has held Florida. Not an election result, just a rumour about his love life... #USElection2016"
kealacove|AltStreamMedia|0.7328|0.0|0.661|0.339|RT @AltStreamMedia: Exit poll favors Trump: Voters most want a 'strong leader' as POTUS https://t.co/Fzk8NDU41N via @MailOnline #Election
kealacove|dailymail|0.7328|0.0|0.661|0.339|RT @AltStreamMedia: Exit poll favors Trump: Voters most want a 'strong leader' as POTUS https://t.co/Fzk8NDU41N via @MailOnline #Election
SWEET_VERGUBA|SWEET_VERGUBA|0.0|0.0|1.0|0.0|"RT @SWEET_VERGUBA: It's finally Election Day! Time to fess up, who are YOU voting for?"
z_jadiazz6|FT|0.0|0.0|1.0|0.0|RT @FT: Latest from @fastFT: Mexican peso climbs further with all eyes on US election https://t.co/cjl6ZrcmxD https://t.co/QX4ImXxP7Y
z_jadiazz6|ft|0.0|0.0|1.0|0.0|RT @FT: Latest from @fastFT: Mexican peso climbs further with all eyes on US election https://t.co/cjl6ZrcmxD https://t.co/QX4ImXxP7Y
BugKlr|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
BugKlr|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
UTnewsie|firstdraftnews|0.4215|0.0|0.882|0.118|"RT @firstdraftnews: If there are stories that made you think ""WOAH"" this election day, take a minute to see if they're true https://t.co/gt"
UTnewsie|t|0.4215|0.0|0.882|0.118|"RT @firstdraftnews: If there are stories that made you think ""WOAH"" this election day, take a minute to see if they're true https://t.co/gt"
SomitraButalia|twitter|0.0|0.0|1.0|0.0|Tune in to KCAL9 news at 4pm for election coverage! https://t.co/1OYYYrXJJy
GreillyPost|CNNnewsroom|0.1027|0.0|0.938|0.063|"RT @CNNnewsroom: The Empire State Building is illuminated in red, white and blue as the candidates await results 1.5 miles apart https://t."
GreillyPost||0.1027|0.0|0.938|0.063|"RT @CNNnewsroom: The Empire State Building is illuminated in red, white and blue as the candidates await results 1.5 miles apart https://t."
AllyJanelle|enoughelise|-0.5106|0.121|0.879|0.0|"RT @enoughelise: if this election has taught me anything, it's that i'm sick of being quiet around my family when it comes to my beliefs."
nadine_morton|smh|0.9169|0.0|0.602|0.398|Great map of the USA showing states won in the race to the White House https://t.co/FhMJVqLru1 #electionday Great map by @smh
nadine_morton|smh|0.9169|0.0|0.602|0.398|Great map of the USA showing states won in the race to the White House https://t.co/FhMJVqLru1 #electionday Great map by @smh
Diggrich_|jpmzo|0.0|0.0|1.0|0.0|RT @jpmzo: Officials: Trump Ballots Switch to Clinton in PA. #VoteFraud. #ElectionFraud. https://t.co/m14QiAgnhR
Diggrich_|breitbart|0.0|0.0|1.0|0.0|RT @jpmzo: Officials: Trump Ballots Switch to Clinton in PA. #VoteFraud. #ElectionFraud. https://t.co/m14QiAgnhR
harobednosyarg|twitter|0.0|0.0|1.0|0.0|"""Grayson, how are you spending your election night?"" https://t.co/y93vQIYXyF"
LessGovt_Now|thefederalistpapers|-0.4019|0.252|0.748|0.0|Voting Machine Error Switching GOP Votes To Democratic https://t.co/pjzdXBToBk
Stepto|synackpse|0.0|0.0|1.0|0.0|@synackpse i think this is the first election it will really show
AlliWriterGirl|recode|0.5423|0.0|0.757|0.243|"People can get free or discounted Uber, Lyft or Zipcar rides to the polls https://t.co/E2Wkv0SSMV https://t.co/fFQ48pqxGU"
carlosgarijo|theverge|0.0|0.0|1.0|0.0|10 provocative political novels to read after the election https://t.co/YrrJoAmppI https://t.co/JyFTsTAjPo
Intashan_C|HuffPostPol|0.0|0.0|1.0|0.0|RT @HuffPostPol: And follow our live analysis right here: https://t.co/PmkRCmLxFx #election https://t.co/7CSTTdsvCp
Intashan_C|huffingtonpost|0.0|0.0|1.0|0.0|RT @HuffPostPol: And follow our live analysis right here: https://t.co/PmkRCmLxFx #election https://t.co/7CSTTdsvCp
ivrosee|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
aydooon|AZegar96|-0.4767|0.185|0.754|0.062|"RT @AZegar96: What's Election Day without an encounter with a racist Trump supporter? Insult me, but just know I'm much more educated than"
FarmerGedon|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
grahampattrsn98|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
manefaemelyano2|reuters|0.0|0.0|1.0|0.0|Reuters: RT ReutersPolitics: Factbox: State-by-state poll closing times for U.S. election https://t.co/u9ISwOiszy https://t.co/Di31h66DTr
KonaTony27|HillaryClinton|0.6114|0.0|0.6|0.4|RT @HillaryClinton: Happy Election Day! https://t.co/jfd3CXLD1s https://t.co/IfOBRuvQzJ
KonaTony27|hillaryclinton|0.6114|0.0|0.6|0.4|RT @HillaryClinton: Happy Election Day! https://t.co/jfd3CXLD1s https://t.co/IfOBRuvQzJ
RobBrimacombe|twitter|0.0|0.0|1.0|0.0|Either way we're gonna need to close one eye and be squeamish!Election all the way. The Canucks have 82. https://t.co/P4wIJxXRSD
JimmyBranley|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
JimmyBranley|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
TarkatanBeauty|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
cumondad|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
cumondad|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
StevenAeons|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
StevenAeons|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
tbishop02|Coop_Engnes2|0.2732|0.0|0.87|0.13|RT @Coop_Engnes2: @natmhef well maybe you'll be old enough to vote in the next election
election_votes|iWafflelicious|0.0|0.0|1.0|0.0|RT @iWafflelicious: Who are you guys voting for?
oweeeneatspears|KdTrey5JR|-0.296|0.104|0.896|0.0|RT @KdTrey5JR: Don't let this election distract you from the fact that the Warriors blew a 3-1 lead in the Finals
SCovitz|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
LocalMarket9|9NEWS|0.2023|0.119|0.714|0.167|RT @9NEWS: Stuck in a line to vote? Here some entertainment while you wait: https://t.co/PQcmFhmWv7
LocalMarket9|9news|0.2023|0.119|0.714|0.167|RT @9NEWS: Stuck in a line to vote? Here some entertainment while you wait: https://t.co/PQcmFhmWv7
envez|cnni|0.0|0.0|1.0|0.0|RT @cnni: Celebrities show off their voting stickers after heading to the polls https://t.co/T98hc03I0a #ElectionNight https://t.co/GIwypoa
envez|cnn|0.0|0.0|1.0|0.0|RT @cnni: Celebrities show off their voting stickers after heading to the polls https://t.co/T98hc03I0a #ElectionNight https://t.co/GIwypoa
mbaangluuc|DonaldJTrumpJr|0.8439|0.062|0.62|0.318|RT @DonaldJTrumpJr: No excuse not to vote. It is your duty to do everything you can to help save America. We can win this thing! #MAGA #Ele
TrumpNewsAlerts|cat_1012000|-0.1531|0.158|0.714|0.128|"RT @cat_1012000: Election Day PrayerLord, We Thank UFor #TrumpPence16Hear our prayer.The wrong shall failThe right prevail#Christians"
rcksk8mech|Jason_Zucker16|0.7755|0.0|0.71|0.29|RT @Jason_Zucker16: Good thing he's better at football than hockey! Don't forget to vote for  @KyleRudolph82 after you vote in today's elec
zagatam|twitter|0.0|0.0|1.0|0.0|Election night Greek food https://t.co/DypSCN0pPJ
Kiko_B7S|YouTube|0.4215|0.0|0.797|0.203|I liked a @YouTube video https://t.co/R0lSqkxdxo The Tale of Election 2016 w/ Benedict Cumberbatch
Kiko_B7S|youtube|0.4215|0.0|0.797|0.203|I liked a @YouTube video https://t.co/R0lSqkxdxo The Tale of Election 2016 w/ Benedict Cumberbatch
alpha_joe86|TeamTrump|0.5574|0.0|0.777|0.223|RT @TeamTrump: 'First Exit Poll: Twice as Many Voters in 2016 Want Strong Leader as President' #ElectionDay https://t.co/pL8TWamWSt
alpha_joe86|breitbart|0.5574|0.0|0.777|0.223|RT @TeamTrump: 'First Exit Poll: Twice as Many Voters in 2016 Want Strong Leader as President' #ElectionDay https://t.co/pL8TWamWSt
BrittanyFlore16|TheChainsmokers|0.0|0.0|1.0|0.0|RT @TheChainsmokers: lets get a little early chainsmoker election poll going... Trump or Hillary... vote below
NathannDH|twitter|-0.1531|0.176|0.682|0.142|This woman on the election news looks like the head from Art Attack https://t.co/32s2HAk74d
DanielleWaldron|postcrescent|0.4199|0.0|0.682|0.318|"Celebrities, they're just like us! #ElectionNight https://t.co/3YzV6ZYpT0"
SiouxCityIow|siouxlandmatters|0.0516|0.0|0.864|0.136|Siouxland Matters Morningside College students bring Sioux City a four hour live Siouxland Matters https://t.co/xDJAEogEtA #SiouxCity #Iowa
ash_atkinson|NickelodeonTV|0.1935|0.158|0.649|0.193|So @NickelodeonTV got super real about election night with their Henry Danger Chip Vote analogy #ElectionNight
12Gage96|Arkansas_Logo|0.0|0.0|1.0|0.0|"RT @Arkansas_Logo: Issue that went unnoticed during this election is how Fayetteville has 80,000 people &amp; only 1 PopeyesCC: @HillaryClinto"
CampSol|instagram|0.6467|0.0|0.72|0.28|We made it! Happy Election Day!  #digital #politics #election2016 #lifeatCS https://t.co/PB7FE5sIr6 https://t.co/i1amaLz2bH
smlyc|JenAshleyWright|0.3612|0.0|0.894|0.106|RT @JenAshleyWright: This election feels like a reminder that the most qualified woman is seen as about as qualified as the least qualified
zumikiss|YasmineGalenorn|0.0|0.0|1.0|0.0|RT @YasmineGalenorn: Our election has now turned deadly. Trump got what he wanted and incited. https://t.co/J0I7bqgzny
zumikiss|twitter|0.0|0.0|1.0|0.0|RT @YasmineGalenorn: Our election has now turned deadly. Trump got what he wanted and incited. https://t.co/J0I7bqgzny
youabu|kickstarter|0.0|0.0|1.0|0.0|Already over the election? I could use your feedback on how my kickstarter page looks. You can preview here:... https://t.co/dD9t8ZI18H
aadair96|jenaeliberty|-0.34|0.156|0.844|0.0|RT @jenaeliberty: I blame my edgy mood on this edgy election #vote2016 #ass #totalass #fuck
DaniloBrack|twitter|0.466|0.0|0.81|0.19|If Democrats like socialism so much...why don't they move to a socialist country???#hypocrisy #election https://t.co/ZMKfc0VqOs
FOX5Vegas|fox5vegas|0.0|0.0|1.0|0.0|Election coverage starts now on #FOX5Vegas &gt;https://t.co/46T2TIPzgX https://t.co/7TTqhO8xHc
BrendaYahm|fox5vegas|0.0|0.0|1.0|0.0|Election coverage starts now on #FOX5Vegas &gt;https://t.co/cp1h0MBWWi https://t.co/XYP3cfPTLa
Trivinho_11|MelissaJoanHart|-0.1531|0.162|0.714|0.123|RT @MelissaJoanHart: Is the election rigged? (Wait for the johnson cameo) ;) https://t.co/AOmf7idEDm
Trivinho_11|twitter|-0.1531|0.162|0.714|0.123|RT @MelissaJoanHart: Is the election rigged? (Wait for the johnson cameo) ;) https://t.co/AOmf7idEDm
Big_Rob2516|BIackPplVids|0.5719|0.0|0.748|0.252|RT @BIackPplVids: Back in 2012 when Obama won the 2012 election  https://t.co/nvEENKBnqj
Big_Rob2516|twitter|0.5719|0.0|0.748|0.252|RT @BIackPplVids: Back in 2012 when Obama won the 2012 election  https://t.co/nvEENKBnqj
jamescass3|MikeDrucker|0.4404|0.0|0.888|0.112|"RT @MikeDrucker: If you have time today, go back and watch some of @LateNightSeth's closer look segments and witness how good he's been thi"
PhonthipC|UberFacts|0.0|0.0|1.0|0.0|RT @UberFacts: Today is Election Day... Take your pick!
RuthHalleran|ForTrump|0.3182|0.0|0.909|0.091|RT @ForTrump: Please get out and vote. Do not listen 2exit polls. This is the election that will decide our country's future.  Let's #MAGA
freeandfunny14|NewsweekEurope|0.0|0.0|1.0|0.0|RT @NewsweekEurope: Read Julian Assange's statement on why Wikileaks has published Clinton campaign documents https://t.co/ojoq2RmEpV https
freeandfunny14|newsweek|0.0|0.0|1.0|0.0|RT @NewsweekEurope: Read Julian Assange's statement on why Wikileaks has published Clinton campaign documents https://t.co/ojoq2RmEpV https
AaronSWillz|HillaryClinton|0.0|0.0|1.0|0.0|Whoever is staying up to watch the US election @HillaryClinton Vs @realDonaldTrump DM me or hmu 
LocalMarket9|9NEWS|0.5411|0.0|0.838|0.162|RT @9NEWS: Enjoy this artist painting the Denver skyline for a moment of zen before election results come in! https://t.co/YINerjIZ1t
LocalMarket9|facebook|0.5411|0.0|0.838|0.162|RT @9NEWS: Enjoy this artist painting the Denver skyline for a moment of zen before election results come in! https://t.co/YINerjIZ1t
MMASOCCERFAN|ananavarro!|0.8016|0.0|0.644|0.356|You're the best thing that came out of Republican party this election cycle ms @ananavarro!
JacqAlex|TheEllenShow|0.4588|0.0|0.857|0.143|"If only Ellen DeGeneres @TheEllenShow was up for election, it would be done and dusted by now. #Election2016 :)"
__Your_Lily|CNNPolitics|-0.2924|0.127|0.873|0.0|"RT @CNNPolitics: On #ElectionDay, Donald Trump still signals he may not accept the results https://t.co/AOUBJX3lqM https://t.co/ngeSYZwbNx"
__Your_Lily|cnn|-0.2924|0.127|0.873|0.0|"RT @CNNPolitics: On #ElectionDay, Donald Trump still signals he may not accept the results https://t.co/AOUBJX3lqM https://t.co/ngeSYZwbNx"
carlgregg|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
Erictrevisan1|mitchellvii|0.5267|0.0|0.848|0.152|"RT @mitchellvii: Democracy Institute, ONLY pollster to correctly guess Brexit, has Trump winning by 5.  Same as my prediction:  https://t.c"
Erictrevisan1||0.5267|0.0|0.848|0.152|"RT @mitchellvii: Democracy Institute, ONLY pollster to correctly guess Brexit, has Trump winning by 5.  Same as my prediction:  https://t.c"
Lonestar357|WordSmithGuy|0.0|0.0|1.0|0.0|RT @WordSmithGuy: Florida Panhandle &amp; Michigan: You have 1 hour &amp; 15 minutes to make history. This entire election may be decided by you gu
justinelturner1|fivethirtyeight|0.4215|0.0|0.865|0.135|"As you start to see how different demographic groups voted this year, it might be helpful to see https://t.co/Dblyqj7WyU"
arruniel|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
arruniel|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
katieli74|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
katieli74|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
deja1422|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
deja1422|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
MikaelaBunker|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: The 15 states that will decide the presidential election https://t.co/SKVjArKSLs https://t.co/rBrxgd8eao
MikaelaBunker|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: The 15 states that will decide the presidential election https://t.co/SKVjArKSLs https://t.co/rBrxgd8eao
lauralong1999|levilusko|0.9209|0.0|0.622|0.378|RT @levilusko: Government positions will always change but the good thing about our great God is:He is never up for re-election. He stands
RockyJeterWebb|KeeganAllen|0.6249|0.0|0.843|0.157|"RT @KeeganAllen: Instead of looking at this election as a series finale of the Great American reality show, look at it as your life...start"
EmilyHug|totalfratmove|0.0|0.0|1.0|0.0|RT @totalfratmove: There is a third option. https://t.co/aNqPlScb9e
EmilyHug|totalfratmove|0.0|0.0|1.0|0.0|RT @totalfratmove: There is a third option. https://t.co/aNqPlScb9e
saharmali|politico|0.2732|0.0|0.811|0.189|Are ya well Kentucky?Trump leads #KYPres; 4.3% reporting. https://t.co/dZ5RN96jca #election2016
freebird_Pepper|Jonbuckhouse|0.6239|0.0|0.843|0.157|RT @Jonbuckhouse: The Polls are starting to close all over the US! Who do you think will win the election?  #ElectionNight #electionday #iV
ThPresident|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
ThPresident|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
efairhurst|youtube|0.0|0.0|1.0|0.0|RNC strategist Sean Spicer offers election night predictions https://t.co/ZYPJaqkO43
nicolemeisner98|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
nicolemeisner98|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
Risefromthedeep|weatherchannel|0.6908|0.0|0.759|0.241|"The @weatherchannel has an ""Escape the Election"" TV music stream rn ""Clouds, rainbows, autumn splendor and smooth jazz evoke tranquility."""
CateStern|twitter|0.0|0.0|1.0|0.0|Watching election results come in tonight https://t.co/TtmSAH6aWc
NathanWalters9|YouTube|0.5319|0.0|0.744|0.256|"Minecraft -(LIVE) ELECTION 2016 ""HELP Build TRUMP'S Wall"": https://t.co/tWckyrSPev via @YouTube"
NathanWalters9|youtube|0.5319|0.0|0.744|0.256|"Minecraft -(LIVE) ELECTION 2016 ""HELP Build TRUMP'S Wall"": https://t.co/tWckyrSPev via @YouTube"
laughingnikki|Capitals|0.0|0.0|1.0|0.0|Im Tweeting to #VoteWilson for @Capitals bobblehead night! Visit https://t.co/8bRp16ujRc for more details! #CapsElectionNight
laughingnikki|nhl|0.0|0.0|1.0|0.0|Im Tweeting to #VoteWilson for @Capitals bobblehead night! Visit https://t.co/8bRp16ujRc for more details! #CapsElectionNight
Hellchick|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
danmccarvel|davidicke|-0.4588|0.176|0.824|0.0|RT @davidicke: This Election Has Disgraced The Entire Profession Of Journalism https://t.co/P0MIuwidcd #Clinton #Trump https://t.co/877waF5
danmccarvel|davidicke|-0.4588|0.176|0.824|0.0|RT @davidicke: This Election Has Disgraced The Entire Profession Of Journalism https://t.co/P0MIuwidcd #Clinton #Trump https://t.co/877waF5
LincolnCleaning|time|-0.4767|0.291|0.709|0.0|"Donald Trump Warns of Voting Problems Nationwide, But Evidence Is Scant https://t.co/6sEtCpeYfA"
gigawell|Stepto|0.5859|0.0|0.833|0.167|@Stepto oddly enough this was my first election season with a land line. Still didn't get polled. I call that a win. Kinda
LRedderso|FredZeppelin12|0.25|0.0|0.895|0.105|RT @FredZeppelin12: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERS. Advantage #Trump. Evening voters are evening voters because t
Robbie_OR|TBNSport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
Robbie_OR|tbnsport|0.2263|0.0|0.899|0.101|RT @TBNSport: Gunnersaurus leapfrogs Clinton and Trump in exit polls as late Arsenal vote proves decisive https://t.co/RddHtb6SxS https://t
desdude_|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
desdude_|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
nicolas_px|becnepla|0.0|0.0|1.0|0.0|RT @becnepla: election news https://t.co/6tk0KK4ZEw
nicolas_px|twitter|0.0|0.0|1.0|0.0|RT @becnepla: election news https://t.co/6tk0KK4ZEw
gaytrashvoid|SICKOFWOLVES|0.0|0.0|1.0|0.0|RT @SICKOFWOLVES: INSTEAD OF HAVING AN ELECTION HAS ANYONE CONSIDERED SPRINTING INTO THE WOODS AND NEVER RETURNING
ShakeYa_Ash|Cartel__shoota|-0.1027|0.119|0.779|0.102|"RT @Cartel__shoota: Waiting on the election results is like waiting for a grade on a group project. I know I did right , I'm scared y'all f"
waltonmolly88|zschwartz11|-0.2263|0.147|0.853|0.0|RT @zschwartz11: They stopped reporting on the election for me. #Blessed https://t.co/pmtnGBwUk3
waltonmolly88|twitter|-0.2263|0.147|0.853|0.0|RT @zschwartz11: They stopped reporting on the election for me. #Blessed https://t.co/pmtnGBwUk3
alden_sia|kolbikay|0.0|0.0|1.0|0.0|". @kolbikay on election day, ""Wait what's a pence?"""
baikal|JonErlichman|0.0|0.0|1.0|0.0|RT @JonErlichman: Things that didn't exist election night in 2008:UberiPadInstagramSnapchatWhatsAppPinterestPeriscopeOculusSlack
RonSpencerRE|realtor|0.6052|0.0|0.78|0.22|Election? What Election?! Check Out These Cute Animals We Found in Listing Photos! https://t.co/trdb6ddGtK https://t.co/B8oWX6oGYK
EnderTheMemelor|barnabybabybump|0.0|0.0|1.0|0.0|RT @barnabybabybump: got my election sticker for tomorrow https://t.co/QQ6myPejGO
EnderTheMemelor|twitter|0.0|0.0|1.0|0.0|RT @barnabybabybump: got my election sticker for tomorrow https://t.co/QQ6myPejGO
manatrue|RT_America|-0.7717|0.34|0.66|0.0|"RT @RT_America: BREAKING: Reports of one dead after gunman opened fire in Azusa, CA https://t.co/G0cuZ0bfH0"
manatrue|rt|-0.7717|0.34|0.66|0.0|"RT @RT_America: BREAKING: Reports of one dead after gunman opened fire in Azusa, CA https://t.co/G0cuZ0bfH0"
bethiecarrillo|twitter|0.0|0.0|1.0|0.0|Election forecast by Tiny https://t.co/wWLbnwSJ2D
infinate_bp|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
Kristi_Craig|G_Eazy|0.7644|0.0|0.752|0.248|"RT @G_Eazy: PLEASE GO OUT AND VOTE WHATEVER YOU DO, THIS COULD BE THE MOST IMPORTANT ELECTION OF OUR LIVES #imwithher #fuckdonaldtrump"
jakobe_luberda|WORLDSTAR|0.5859|0.0|0.678|0.322|RT @WORLDSTAR: Who will win the 2016 presidential election? 
slvrfnx|ABC|0.0|0.0|1.0|0.0|RT @ABC: ELECTION NIGHT: Who will be our next president? Coverage starting at 7PM ET on @ABCNetwork and across @ABC digital: https://t.co/V
slvrfnx|t|0.0|0.0|1.0|0.0|RT @ABC: ELECTION NIGHT: Who will be our next president? Coverage starting at 7PM ET on @ABCNetwork and across @ABC digital: https://t.co/V
JohnnyTruax|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
DAnnRenn|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
DAnnRenn||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
jhallang|ABC|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
jhallang|abcnews|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
manefaemelyano2|reuters|0.0|0.0|1.0|0.0|Reuters: RT ReutersPolitics: Former President George W. Bush does not cast vote for president https://t.co/pZNdPY7GeP
Chance_Takers|twitter|0.2225|0.0|0.914|0.086|We're back on FB Live! Want to know the second weed gets legalized? IGH TIMES is covering the election live! https://t.co/dCB4oHO97v
RickMitchellWX|twitter|0.0|0.0|1.0|0.0|Fueling up for a busy night of election coverage. #nbcdfw https://t.co/fRok4sVbsN
the_gxdess|abiriketaa|0.8074|0.0|0.733|0.267|"RT @abiriketaa: Every time I think I of Donald trump winning the election I hear ""blessed be our new founding fathers for letting us purge."
jorgee3169|STXR67|0.4767|0.0|0.871|0.129|RT @STXR67: RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exc
CodyPhelan|FT|0.0|0.0|1.0|0.0|RT @FT: It's Trump vs Clinton: how did the US election polls end up? https://t.co/Ih7NEPtbfK https://t.co/7WxqAO4IWS
CodyPhelan|ig|0.0|0.0|1.0|0.0|RT @FT: It's Trump vs Clinton: how did the US election polls end up? https://t.co/Ih7NEPtbfK https://t.co/7WxqAO4IWS
garethjhill|garethjhill|-0.1546|0.182|0.682|0.136|Silliest election ever? And not in a good way. https://t.co/CClR8aIq8Y #ElectionNight https://t.co/3BJkqhtFrI
SamnangMedia|ABCNews24|0.4404|0.0|0.861|0.139|RT @ABCNews24: Will the sleeping giant wake &amp; change this election? @chas_usa discusses the influential latino vote #usavotes https://t.co/
SamnangMedia|t|0.4404|0.0|0.861|0.139|RT @ABCNews24: Will the sleeping giant wake &amp; change this election? @chas_usa discusses the influential latino vote #usavotes https://t.co/
Arlhet_Stranger|AllyBrooke|0.7506|0.0|0.575|0.425|RT @AllyBrooke: Praying for our election tomorrow and may God bless our country 
3Dstoretn|3dprint|0.0|0.0|1.0|0.0|3Dstore.tn US Election 2016: The Washington Post to 3D Print Results Live https://t.co/CwYXi5m6dB https://t.co/WKbIXqALvl
kysgabbygirl|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
InTheSoupAgain|BBCRadio4|0.7772|0.0|0.625|0.375|"Listening to @BBCRadio4 election new special. Rather good, not as depressing as I thought it would be."
travisbernard|twitter|0.4939|0.0|0.714|0.286|This cant be rightelection coverage looks pretty tasty. https://t.co/qB6fjqLL2O
peacematters2|Verge|0.0516|0.242|0.466|0.292|"Want a good, healthy cry? Watch the live stream of Susan B. Anthonys grave https://t.co/aMXCp67ZOL via @Verge"
peacematters2|theverge|0.0516|0.242|0.466|0.292|"Want a good, healthy cry? Watch the live stream of Susan B. Anthonys grave https://t.co/aMXCp67ZOL via @Verge"
1913Facts|Chicagoist|0.1027|0.103|0.769|0.128|RT @Chicagoist: Chicago Remembers Suffragist Badass Ida B. Wells On Election Day https://t.co/YyRAbcSqNt https://t.co/yopczX8sho
1913Facts|chicagoist|0.1027|0.103|0.769|0.128|RT @Chicagoist: Chicago Remembers Suffragist Badass Ida B. Wells On Election Day https://t.co/YyRAbcSqNt https://t.co/yopczX8sho
ThatDickScott|john_wawrow|-0.2411|0.179|0.821|0.0|@john_wawrow I'm not sure he's a part of election night coverage.
kjb568|voguemagazine|0.0|0.0|1.0|0.0|RT @voguemagazine: We're #withher. https://t.co/MaeV79cEhz https://t.co/wsWRxIAdxq
kjb568|vogue|0.0|0.0|1.0|0.0|RT @voguemagazine: We're #withher. https://t.co/MaeV79cEhz https://t.co/wsWRxIAdxq
8_christiansen|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
jbonner49|PaperWash|0.3612|0.0|0.878|0.122|RT @PaperWash: Here is what the electoral map would look like if only millennials voted in the election https://t.co/QSialAhyEx
jbonner49|twitter|0.3612|0.0|0.878|0.122|RT @PaperWash: Here is what the electoral map would look like if only millennials voted in the election https://t.co/QSialAhyEx
Auttiee_|robbins_dexter|-0.4574|0.207|0.655|0.138|RT @robbins_dexter: No matter the result of the election or how good or bad things get Jesus Christ is still on the throne! 
Byone028|NorahODonnell|0.0|0.0|1.0|0.0|"RT @NorahODonnell: After 18 months, were finally here, Election Night 2016, tune into our coverage (7PM ET): https://t.co/wTIcGIzmeE!"
Byone028|cbsnews|0.0|0.0|1.0|0.0|"RT @NorahODonnell: After 18 months, were finally here, Election Night 2016, tune into our coverage (7PM ET): https://t.co/wTIcGIzmeE!"
hannahyonks|Things4WhitePpl|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
hannahyonks|twitter|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
cwsparker|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
cwsparker|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
DeAngelisNews|washingtonpost|0.0|0.0|1.0|0.0|News: Donald Trump was booed before he voted for Donald Trump - Washington Post https://t.co/qFPfElmDoc
Gww1863|geekybeergal|0.8478|0.0|0.566|0.434|RT @geekybeergal: Happy Election Day! I can pretty much guarantee we'll all be drinking tonight. https://t.co/9cykNFoQk6
Gww1863|facebook|0.8478|0.0|0.566|0.434|RT @geekybeergal: Happy Election Day! I can pretty much guarantee we'll all be drinking tonight. https://t.co/9cykNFoQk6
Dr_C2006|mamapojo|0.8834|0.0|0.671|0.329|"RT @mamapojo: Watching early election results: If HRC wins I'll go to bed, sleep better; if DT wins I finish this bottle while googling hou"
brire04|JoeyGraceffa|0.5461|0.0|0.773|0.227|RT @JoeyGraceffa: RT IF YOU'RE READY FOR THIS ELECTION TO BE OVER!  #ImWithHer
YoursTrulyHer0|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
YoursTrulyHer0|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
jashwat07|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
jashwat07|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
Ddebn8R|markos|-0.0572|0.067|0.933|0.0|"RT @markos: CNN exit poll, 38% wanted change. That's not the number Trump needed. This wasn't a change election."
Thejeepboss|ashlynbradnerr|0.0|0.0|1.0|0.0|"RT @ashlynbradnerr: enough about the election, look at the jeep  https://t.co/Sa2ZFsvfQi"
Thejeepboss|twitter|0.0|0.0|1.0|0.0|"RT @ashlynbradnerr: enough about the election, look at the jeep  https://t.co/Sa2ZFsvfQi"
CamaroKiddos|DonaldJTrumpJr|0.4753|0.0|0.894|0.106|RT @DonaldJTrumpJr: The easiest way to get my father to do something is tell him it can't be done! Today we take back America from the elit
jenthegoat|_elsti_|-0.4341|0.207|0.793|0.0|RT @_elsti_: I have never been so worried about politics until this election
marytg66|UpshotNYT|0.5859|0.0|0.725|0.275|RT @UpshotNYT: When will we know we have a winner? https://t.co/1pMJXK7mS4 https://t.co/B87hwbBQZy
marytg66|nytimes|0.5859|0.0|0.725|0.275|RT @UpshotNYT: When will we know we have a winner? https://t.co/1pMJXK7mS4 https://t.co/B87hwbBQZy
efairhurst|mashable|0.0|0.0|1.0|0.0|America gets lit: The Lite Brite guide to election results https://t.co/KOXFQJ3LLx
itsleovalentino|YouTube|0.4215|0.0|0.797|0.203|I liked a @YouTube video https://t.co/jZIjx6txyF Decision 2016: LIVE Election Night Coverage | NBC News
itsleovalentino|youtube|0.4215|0.0|0.797|0.203|I liked a @YouTube video https://t.co/jZIjx6txyF Decision 2016: LIVE Election Night Coverage | NBC News
Jean0x|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
bherbst33|CTVVancouver|0.4019|0.0|0.787|0.213|RT @CTVVancouver: LIVE @ 4 p.m.: America's Choice 2016 election special. https://t.co/ygNE6FxwXa https://t.co/QNZ5P7bG3O
bherbst33|bc|0.4019|0.0|0.787|0.213|RT @CTVVancouver: LIVE @ 4 p.m.: America's Choice 2016 election special. https://t.co/ygNE6FxwXa https://t.co/QNZ5P7bG3O
_succ_papi_|Drops|0.6633|0.0|0.793|0.207|RT @Drops: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  LOS ANGELES
JSCram3254|jonrog1|0.8395|0.0|0.68|0.32|RT @jonrog1: The most adorable way to track - love the County profiles when you zoom in!  https://t.co/SIvBetE3V6 via @GuardianUS
JSCram3254|theguardian|0.8395|0.0|0.68|0.32|RT @jonrog1: The most adorable way to track - love the County profiles when you zoom in!  https://t.co/SIvBetE3V6 via @GuardianUS
2k_joseph|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
2k_joseph|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
davegisaac|JasonAlt_dj|0.0|0.0|1.0|0.0|"RT @JasonAlt_dj: ELECTION 2016: Your one-stop place for results from Camden, Burlington &amp; Gloucester counties https://t.co/Zx5z0zEba0"
davegisaac|courierpostonline|0.0|0.0|1.0|0.0|"RT @JasonAlt_dj: ELECTION 2016: Your one-stop place for results from Camden, Burlington &amp; Gloucester counties https://t.co/Zx5z0zEba0"
JeffMcClelland|alyankovic|0.5312|0.0|0.847|0.153|"RT @alyankovic: What, it's Election Day ALREADY?? Man, that campaign season just FLEW BY!!!!!! Okay, America, let's do this. https://t.co/t"
JeffMcClelland|twitter|0.5312|0.0|0.847|0.153|"RT @alyankovic: What, it's Election Day ALREADY?? Man, that campaign season just FLEW BY!!!!!! Okay, America, let's do this. https://t.co/t"
OmarjSakr|twitter|0.5267|0.115|0.635|0.25|"Take a break from election madness, read a poem. A poem about family, love, boys, god &amp; country. How they rupture. https://t.co/bqRaAntHYr"
xo_leahbrown_xo|GavinReacts|0.6249|0.0|0.661|0.339|RT @GavinReacts: A great way to start Election Day https://t.co/OWJDlMLbs5
xo_leahbrown_xo|twitter|0.6249|0.0|0.661|0.339|RT @GavinReacts: A great way to start Election Day https://t.co/OWJDlMLbs5
diawrites|YouTube|0.0|0.0|1.0|0.0|Decision 2016: LIVE Election Night Coverage | NBC News https://t.co/nI4xp7C5IW via @YouTube
diawrites|youtube|0.0|0.0|1.0|0.0|Decision 2016: LIVE Election Night Coverage | NBC News https://t.co/nI4xp7C5IW via @YouTube
ScottFralick|BoyerMichel|0.0|0.0|1.0|0.0|RT @BoyerMichel: CTV Edmonton election coverage from the Garneau theatre tonight! Live in just a few! @ctvedmonton https://t.co/NTTm5qvU4x
ScottFralick|twitter|0.0|0.0|1.0|0.0|RT @BoyerMichel: CTV Edmonton election coverage from the Garneau theatre tonight! Live in just a few! @ctvedmonton https://t.co/NTTm5qvU4x
CarinaNicole16|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
CarinaNicole16|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
alexn_leigh|JustinWolfers|0.6908|0.0|0.749|0.251|"RT @JustinWolfers: By the power vested in me by F**kface Von Clownstick, I hereby declare it a special Election Day beer o'clock for the ha"
debbiedo58|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
xoxotabello|ddlovato|0.1027|0.101|0.734|0.165|RT @ddlovato: I apologize for the joke I made earlier.. seemed to offend some people. Just making light of the election 
sophie_js|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
sophie_js|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
Nathalielassus1|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: The latest updates on the House races https://t.co/Q1iwJbI6El https://t.co/SvkRA88ctf
Nathalielassus1|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: The latest updates on the House races https://t.co/Q1iwJbI6El https://t.co/SvkRA88ctf
Margie_Burns|GOP|0.7717|0.0|0.705|0.295|@GOP https://t.co/Y1lYF63i5A Keep polls open in NC. But not out of false hope that Clinton will win there.
Margie_Burns|margieburns|0.7717|0.0|0.705|0.295|@GOP https://t.co/Y1lYF63i5A Keep polls open in NC. But not out of false hope that Clinton will win there.
syaldram|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
titi_jennie|USATODAY|0.0|0.0|1.0|0.0|RT @USATODAY: 49ers quarterback Colin Kaepernick has chosen to stay on the sidelines for this presidential election. #ElectionNight https:/
titi_jennie||0.0|0.0|1.0|0.0|RT @USATODAY: 49ers quarterback Colin Kaepernick has chosen to stay on the sidelines for this presidential election. #ElectionNight https:/
jdprose|anna_orso|0.3612|0.0|0.865|0.135|RT @anna_orso: Toomey told voters he supports Donald Trump... one hour before polls close in Pennsylvania. https://t.co/l5iThHjOMR
jdprose|billypenn|0.3612|0.0|0.865|0.135|RT @anna_orso: Toomey told voters he supports Donald Trump... one hour before polls close in Pennsylvania. https://t.co/l5iThHjOMR
DanBennett|bbcthree|0.6593|0.0|0.779|0.221|I mean. I get why. But also it's not our election. This would be great on @bbcthree if they didn't screw that up
DomminickG|FunnyPicsDepot|0.0|0.0|1.0|0.0|RT @FunnyPicsDepot: How to start off Election Day right https://t.co/RANxmEYi64
DomminickG|twitter|0.0|0.0|1.0|0.0|RT @FunnyPicsDepot: How to start off Election Day right https://t.co/RANxmEYi64
viralwomen|mic|0.0|0.0|1.0|0.0|Here's when we can expect to learn who the next president will be. Mic https://t.co/fJFhTTkhkX
gocoo|AustinMahone|0.6114|0.0|0.501|0.499|RT @AustinMahone: Happy Election Day! 
scooter_annie|williamderraugh|0.8608|0.0|0.701|0.299|RT @williamderraugh: IF YOU'RE IN FLORIDA AND YOU SUPPORT TRUMP'S AMERICA FIRST POLICIES YOU CAN WIN THIS ELECTION FOR AMERICA! MUST VOTE!
steelcitydavid|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
steelcitydavid|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
andiius_|KathleenLights1|0.4199|0.141|0.573|0.286|RT @KathleenLights1: Hope everyone voted today! This election has traumatized me.... I pray for America.
swankerella|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
swankerella|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
2_3ZoneCoach|bobfescoe|0.0|0.0|1.0|0.0|RT @bobfescoe: So do they know the results of the election in London already?
ColleyKellerCt|CBSDFW|-0.5267|0.167|0.833|0.0|RT @CBSDFW: Dallas County election judge assaulted and robbed Monday night.  Can't work polling place on #ElectionDay. https://t.co/ML8HrAS
ColleyKellerCt|t|-0.5267|0.167|0.833|0.0|RT @CBSDFW: Dallas County election judge assaulted and robbed Monday night.  Can't work polling place on #ElectionDay. https://t.co/ML8HrAS
m_gordon_umc|twitter|0.0|0.0|1.0|0.0|Election night pizza! https://t.co/hEBiFqhSYw
AngelSanchezGDL|LosinDonald|-0.5574|0.247|0.753|0.0|"RT @LosinDonald: Trump distorts CNN report, incorrectly tweets nationwide election results are suspect by @jeisrael https://t.co/wd8sUFbU"
AngelSanchezGDL|t|-0.5574|0.247|0.753|0.0|"RT @LosinDonald: Trump distorts CNN report, incorrectly tweets nationwide election results are suspect by @jeisrael https://t.co/wd8sUFbU"
mhmhart|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
mhmhart||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
IlladelphAC|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
IlladelphAC|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
RobaelEnyew|twitter|0.0|0.0|1.0|0.0|This was at my voting precinct today. Had nothing to do with the election but I realllly wanna know what event this https://t.co/vRpVbm6MEK
ELIZABETHMALTE2|mypchurch|0.5473|0.0|0.694|0.306|RT @mypchurch: ELECTIONRESULTSTONIGHTWe watch as a UNITED NATIONDr Michael Chitwoodhttps://t.co/unyOZJe1
Richnavin86|brookeperrin|0.6876|0.054|0.707|0.239|RT @brookeperrin: I'm so happy about meeting @MarnieTheDog that this election doesn't even matter anymore https://t.co/Bj58Dx3DgE
Richnavin86|twitter|0.6876|0.054|0.707|0.239|RT @brookeperrin: I'm so happy about meeting @MarnieTheDog that this election doesn't even matter anymore https://t.co/Bj58Dx3DgE
ChrisOchsnerKC|KCStarShane|0.0|0.0|1.0|0.0|RT @KCStarShane: Clay Countys District 17 possibly had the longest wait to vote in Kansas City #ElectionDay @KCStar https://t.co/I2IBdAqqt
ChrisOchsnerKC|t|0.0|0.0|1.0|0.0|RT @KCStarShane: Clay Countys District 17 possibly had the longest wait to vote in Kansas City #ElectionDay @KCStar https://t.co/I2IBdAqqt
haleybug741|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
Mariahpatrice__|lorenlondin|-0.4404|0.326|0.674|0.0|RT @lorenlondin: I'm scared about this election 
SpeakYOURmindT|ABCWorldNews|-0.0258|0.096|0.812|0.092|RT @ABCWorldNews: Scores of people are waiting in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.
SpeakYOURmindT||-0.0258|0.096|0.812|0.092|RT @ABCWorldNews: Scores of people are waiting in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.
JWPrairieDog|tulsaworld|0.3818|0.0|0.88|0.12|"Long live #newsroompizza on election nights. As the pizza goes, so goes the newspaper industry. @tulsaworld keeping the tradition alive."
MikeDeVillaer|DemiNewell|0.168|0.0|0.9|0.1|"RT @DemiNewell: ""Do you want to turn on the election coverage?""""Why? It isn't real.""""Good point."" #ElectionNight"
RahsaanBall|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
RahsaanBall|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
JustinGorify|CNN|-0.1531|0.071|0.929|0.0|RT @CNN: Time is running out for @HillaryClinton &amp; @realDonaldTrump. Its a close race. Dont miss a moment on election night with CNN. htt
brenna1009|chelliet22|-0.0772|0.058|0.942|0.0|"RT @chelliet22: ""We're sorry for everything you've had to endure and learn leading up to this election.""Americans, to the world. And ours"
JoeyHopalong|byrdinator|0.0|0.0|1.0|0.0|RT @byrdinator: picking up some refreshments for election night!!! https://t.co/yAaHCOuWey
JoeyHopalong|twitter|0.0|0.0|1.0|0.0|RT @byrdinator: picking up some refreshments for election night!!! https://t.co/yAaHCOuWey
vostokintheair|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
vostokintheair|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
zoe_nor|latimes|0.0|0.0|1.0|0.0|Former President George W. Bush didn't vote for Donald Trump https://t.co/VD14r8IOqb
4Wrath|dissonance_pod|0.0|0.0|1.0|0.0|Are you watching @dissonance_pod 's live coverage of the election?Well you should be: https://t.co/1bDKCXgOZP ~ A
4Wrath|youtube|0.0|0.0|1.0|0.0|Are you watching @dissonance_pod 's live coverage of the election?Well you should be: https://t.co/1bDKCXgOZP ~ A
WillRowland7|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
nhaatt|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
nhaatt|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
DrPepperJutsu|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
DrPepperJutsu|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
TenderThomas|FiveThirtyEight|0.0|0.0|1.0|0.0|RT @FiveThirtyEight: Remember when ... https://t.co/bmwTj0VQYX https://t.co/ViSCxeRhJW
TenderThomas|fivethirtyeight|0.0|0.0|1.0|0.0|RT @FiveThirtyEight: Remember when ... https://t.co/bmwTj0VQYX https://t.co/ViSCxeRhJW
ChipotleGetsMe|dissonance_pod|0.0|0.0|1.0|0.0|RT @dissonance_pod: Watch us watch election TV and stuff: https://t.co/KmED4IDnsk
ChipotleGetsMe|youtube|0.0|0.0|1.0|0.0|RT @dissonance_pod: Watch us watch election TV and stuff: https://t.co/KmED4IDnsk
leria__v|Auburnnn14|0.128|0.14|0.699|0.162|RT @Auburnnn14: Idc who wins the election cuz at the end of the day we screwed ether way
Rich_Laudermilk|ABC|0.0|0.0|1.0|0.0|RT @ABC: ELECTION NIGHT: Who will be our next president? Coverage starting at 7PM ET on @ABCNetwork and across @ABC digital: https://t.co/V
Rich_Laudermilk|t|0.0|0.0|1.0|0.0|RT @ABC: ELECTION NIGHT: Who will be our next president? Coverage starting at 7PM ET on @ABCNetwork and across @ABC digital: https://t.co/V
MicheleJawando|newsone!|0.0|0.0|1.0|0.0|3 minutes until we are live for election night coverage here in DC on @newsone! https://t.co/QQ7wJsMKKE
MicheleJawando|twitter|0.0|0.0|1.0|0.0|3 minutes until we are live for election night coverage here in DC on @newsone! https://t.co/QQ7wJsMKKE
WhoareyouBO|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
Duncks|instagram|0.3612|0.0|0.815|0.185|I'm ready to watch the election results. #wonderwoman #lularoe #imwithher #electionday https://t.co/4ik2Sm1hGL
crowjane29|pastemagazine|0.34|0.0|0.862|0.138|"Samantha Bee Endorses Hillary, Reads Emails and Goes to Russia In Last Pre-Election Full Frontal https://t.co/NXaTAibi8G"
WSBT|wsbt|-0.4019|0.278|0.722|0.0|Live video from battleground state of Ohio: https://t.co/qvdABMlNWV
yjsTm1YVRUupi5j|WDFx2EU8|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
yjsTm1YVRUupi5j|t|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
amishabarnes2|chungaah|0.3818|0.122|0.667|0.211|RT @chungaah: Not even worried about the election Ik who gonna win Hillary obviously 
monseans|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
monseans|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
LG_Noojoya|twitter|0.0|0.0|1.0|0.0|Let the election results begin https://t.co/c4GYgxVonP
goodbyetoyou|GMA|0.0|0.0|1.0|0.0|RT @GMA: MINUTES AWAY: #ElectionNight from Times Square: https://t.co/9FrLR8ogNb https://t.co/A24qjFfpYD
goodbyetoyou|abcnews|0.0|0.0|1.0|0.0|RT @GMA: MINUTES AWAY: #ElectionNight from Times Square: https://t.co/9FrLR8ogNb https://t.co/A24qjFfpYD
nattsurf|twitter|0.5574|0.0|0.783|0.217|These are the funniest memes of the US Election so far - The Sun https://t.co/XLgiJsvlyv
morethanasong5|secure|0.0|0.0|1.0|0.0|"Donald J. Trump for President, Inc. https://t.co/5ilMv8fRIY"
Kress_Golfnut|politico|0.6249|0.0|0.549|0.451|Great site to follow election on:https://t.co/1oJvqotg1d
UrFaceCrunchy|Mr_Spacely_87|0.5859|0.087|0.705|0.208|RT @Mr_Spacely_87: Even tho I'm going the vote.. y'all do kno there has been presidents that won the popular vote and still lose the electi
Kaytaroo|corshit|0.0|0.0|1.0|0.0|@corshit I don't have my phone I'm on Morgan's &amp; we are at my grandparents watching the election
ohmyzan|hyunascult|-0.5214|0.2|0.698|0.103|"@hyunascult like this entire election, even when BERNIE was running, she was all for Hillary so wtf is this"
bettyssd|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Obama continues Election Day ritual for Hillary Clinton https://t.co/uxU8EZ7jC3
bettyssd|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Obama continues Election Day ritual for Hillary Clinton https://t.co/uxU8EZ7jC3
_josie98|AyannaImani13|0.0258|0.151|0.653|0.196|RT @AyannaImani13: I hate radical Christians who act like they weren't having sex earlier today. Go pray over this election. 
_theangellica|dj_rocklee|0.5374|0.082|0.752|0.166|RT @dj_rocklee: Shiiitttt if Donald Trump wins this election im warning ALL YALL !!!!! Knuck if you buck white America. Knuck if you the
danielmarans|EricMarkowitz|0.0|0.0|1.0|0.0|RT @EricMarkowitz: It's the yule log for election night! https://t.co/EeSU8DCTp0
danielmarans|twitter|0.0|0.0|1.0|0.0|RT @EricMarkowitz: It's the yule log for election night! https://t.co/EeSU8DCTp0
TrumpManDoo|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
TrumpManDoo||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
BMacvay|CrystalMoon214|0.0|0.0|1.0|0.0|RT @CrystalMoon214: Watching election coverage like... https://t.co/mE2zW7nQ7A
BMacvay|twitter|0.0|0.0|1.0|0.0|RT @CrystalMoon214: Watching election coverage like... https://t.co/mE2zW7nQ7A
MetteSAndersen|StephenMcGann|0.6249|0.0|0.797|0.203|"RT @StephenMcGann: Never mind the election, here's a nice picture of a badger in my garden, captured on my infra-red night camera :-) https"
devin_ray49|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
JayXombie|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
JayXombie|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
JakeM_1998|twitter|0.0|0.0|1.0|0.0|Stand by for #CNNElection projectionhttps://t.co/4FQCP7mZzp#ElectionNight https://t.co/RTU44TAgpc
NoshFoodandWine|nytimes|0.0|0.0|1.0|0.0|"The Unpublished Poems of Donald J. Trump, 2015-16 https://t.co/weGaCS4pvW"
DianeNC|mitchellvii|0.0|0.0|1.0|0.0|"@mitchellvii Donald Trump Election Night Speech in New York, NY https://t.co/F8HtH0VG0e"
DianeNC|lifezette|0.0|0.0|1.0|0.0|"@mitchellvii Donald Trump Election Night Speech in New York, NY https://t.co/F8HtH0VG0e"
wildwestwalker2|NZStuff|-0.7096|0.312|0.688|0.0|"RT @NZStuff: US election: Shots fired near California polling station, four victims reported https://t.co/kig7RAB6QM https://t.co/Kkai7oIlxO"
wildwestwalker2|stuff|-0.7096|0.312|0.688|0.0|"RT @NZStuff: US election: Shots fired near California polling station, four victims reported https://t.co/kig7RAB6QM https://t.co/Kkai7oIlxO"
StarSuperKai|twitch|-0.5242|0.195|0.805|0.0|LIVE! Continuing Dishonored!Come hang out and chill while you stress about the election &lt;3 https://t.co/hcTp5ntWE2
lindsaytupy|ALLIEineed2P|0.4215|0.092|0.734|0.174|RT @ALLIEineed2P: stuck between wanting the election to be over and not wanting to know the result :-))
svizzman|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
joshuamcgee0325|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
joshuamcgee0325|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
VeeFrancine|RaunchyBillups|-0.296|0.095|0.905|0.0|RT @RaunchyBillups: Can I distract y'all from the election real quick and inform you that Apple Music is indeed for the culture https://t.c
VeeFrancine||-0.296|0.095|0.905|0.0|RT @RaunchyBillups: Can I distract y'all from the election real quick and inform you that Apple Music is indeed for the culture https://t.c
redlyn68|ananavarro|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
redlyn68|twitter|0.0|0.0|1.0|0.0|RT @ananavarro: So I bought a white pantsuit for election coverage tonight about a month ago...before I knew it was a thing. https://t.co/D
zoe_nor|latimes|0.0|0.0|1.0|0.0|How this election has revealed workplace sexism is still an issue https://t.co/FxSOorFMRT
dstys167|Bipartisanism|0.8415|0.0|0.635|0.365|RT @Bipartisanism: Women Do Something AWESOME To Honor Susan B. Anthony On Election Day(DETAILS) https://t.co/WkO2qMGZpd https://t.co/p8xM
dstys167|bipartisanreport|0.8415|0.0|0.635|0.365|RT @Bipartisanism: Women Do Something AWESOME To Honor Susan B. Anthony On Election Day(DETAILS) https://t.co/WkO2qMGZpd https://t.co/p8xM
denlogue|weatherchannel|0.8225|0.0|0.397|0.603|Election night winner? @weatherchannel #EscapetheElection.  Brilliant #fb
backFickle|MVxrse|0.3612|0.0|0.848|0.152|RT @MVxrse: People who really know about the election what's it looking like right now
PrometheusLaw|foreignpolicy|0.7269|0.0|0.664|0.336|ForeignPolicy: RT FPMediaDept: Join djrothkopf NYCComedyCellar &amp; a host of smart &amp; informed media &amp; comedians toni https://t.co/gNDHjlXluX
unlsweetie|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
unlsweetie|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
BrittyDiFitty1|BuzzFeedNews|0.0|0.0|1.0|0.0|"RT @BuzzFeedNews: So far today, there have been 25 million tweets about the election sent through 6pm EST #Election2016"
mowser1970|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
JakeM_1998|snappytv|0.743|0.105|0.576|0.319|"RT AC360: .ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Tr https://t.co/VXcIce2zNV"
SpannaGattinara|joshtpm|0.0|0.0|1.0|0.0|RT @joshtpm: Last time we let Utah run the nationwide election https://t.co/h0bQzw8tMa
SpannaGattinara|twitter|0.0|0.0|1.0|0.0|RT @joshtpm: Last time we let Utah run the nationwide election https://t.co/h0bQzw8tMa
scottu|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
scottu|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
rory_svw|_alastair|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
rory_svw|t|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
carstarr6|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: There have been 25 million tweets sent around the world about the US election today, per @twitter https://t.co/dcOvqM"
carstarr6|t|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: There have been 25 million tweets sent around the world about the US election today, per @twitter https://t.co/dcOvqM"
PablodelaMac|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
PablodelaMac|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
So_Officiial|khendoll|0.0|0.0|1.0|0.0|RT @khendoll: Me waiting for these election results cause I know Twitter about to be popping all night #ElectionNight https://t.co/kOzyUcIE
So_Officiial|t|0.0|0.0|1.0|0.0|RT @khendoll: Me waiting for these election results cause I know Twitter about to be popping all night #ElectionNight https://t.co/kOzyUcIE
rjpanetti|voxdotcom|0.0|0.0|1.0|0.0|RT @voxdotcom: These early states could give us clues about how the rest of the night will go. https://t.co/6MhzzHQKnM https://t.co/NzavKRd
rjpanetti|vox|0.0|0.0|1.0|0.0|RT @voxdotcom: These early states could give us clues about how the rest of the night will go. https://t.co/6MhzzHQKnM https://t.co/NzavKRd
Walk_Like_MoDel|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
jessicabanov|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
jessicabanov|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
miflorhermosa|SInow|0.0|0.0|1.0|0.0|RT @SInow: Colin Kaepernick said he isnt voting in the election https://t.co/9IfZWrKNCc https://t.co/l3kO9BORir
miflorhermosa|si|0.0|0.0|1.0|0.0|RT @SInow: Colin Kaepernick said he isnt voting in the election https://t.co/9IfZWrKNCc https://t.co/l3kO9BORir
Gus_Tinajero4|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
Gus_Tinajero4|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
Moeezus|SirachAbebe|-0.8074|0.399|0.601|0.0|RT @SirachAbebe: This election is sadder than Bing Bong's death in Inside Out
JesseJaymz|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
swann_combs|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
dailydot|dailydot|0.296|0.0|0.804|0.196|"Surviving 2016: Live election results, memes, and news: https://t.co/8Q2q2yU9LY https://t.co/CxX2Ml1bMc"
JSYK|twitter|0.0|0.0|1.0|0.0|"Remember yesterday when i was all ""if only the election were on a non-work day and we could watch election tv all d https://t.co/1tkLQRXBsK"
torisuemagoo|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
torisuemagoo|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
__thatgirlmya|Dex_Jay|0.0|0.0|1.0|0.0|RT @Dex_Jay: Steve Harvey Should Announce The Election 
rynkinazywo|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
rynkinazywo|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
OneLastMyth|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
seniaabeniaa|_ummkeesh|-0.5032|0.146|0.854|0.0|RT @_ummkeesh: Some people are so fucking ignorant about this presidential election! Stfu! educate yourself before you speak on it.
dotlayer8|dailydot|0.296|0.0|0.804|0.196|"Surviving 2016: Live election results, memes, and news: https://t.co/2FbMDtlYqa https://t.co/HcLP2wTgLm"
SculptNewYork|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
MinallSan|JessieJaneDuff|-0.4574|0.125|0.875|0.0|RT @JessieJaneDuff: Volunteers take thousands of Amish voters to the polls in battleground Ohio &amp; PA for a Trump barn raiser! #VoteTrump ht
bwild76|ronnieruff|-0.1531|0.133|0.758|0.11|RT @ronnieruff: Who is going to get high as fuck for Election Night? It will be far better I think  #ElectionNight #ElectionDay #LegalizeCA
YoungCreateers|TheEllenShow|0.0|0.0|1.0|0.0|"@TheEllenShow ""I imagined I voted""!@YoungCreateers #animals #dog #dogs #pet #kids #books #parents #vote https://t.co/NDyTBDqIQA"
YoungCreateers|twitter|0.0|0.0|1.0|0.0|"@TheEllenShow ""I imagined I voted""!@YoungCreateers #animals #dog #dogs #pet #kids #books #parents #vote https://t.co/NDyTBDqIQA"
DebraDianeParr|vivelafra|0.6884|0.0|0.794|0.206|"RT @vivelafra: THE MONSTER VOTE IS REAL!!! &gt;&gt;&gt; Trump Could Win Michigan, Turnout 'Much Higher than Expected' https://t.co/fY1Ex7V8Ot #Trump"
DebraDianeParr|breitbart|0.6884|0.0|0.794|0.206|"RT @vivelafra: THE MONSTER VOTE IS REAL!!! &gt;&gt;&gt; Trump Could Win Michigan, Turnout 'Much Higher than Expected' https://t.co/fY1Ex7V8Ot #Trump"
onlyjustginger|nataliemjb|-0.3595|0.151|0.849|0.0|"RT @nataliemjb: Get your election results here! (No models, no extraneous data, just results) https://t.co/oaJGzR9GeJ"
onlyjustginger|elections|-0.3595|0.151|0.849|0.0|"RT @nataliemjb: Get your election results here! (No models, no extraneous data, just results) https://t.co/oaJGzR9GeJ"
libertad717|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
libertad717|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
DoveyFL|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
DoveyFL||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
mjohnson_music|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
mjohnson_music|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
epitygxanwn|_eric_alexander|-0.4215|0.149|0.851|0.0|"@_eric_alexander Speaking of him, reading 'nausea' upside down, I told pharmacist I thought election atmosphere duped me 2 read 'nutcase'"
Liiids|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Liiids|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
JHoff2214|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
JHoff2214|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
forBittenpeach|suttonimpaQt|0.3612|0.0|0.828|0.172|RT @suttonimpaQt: This election is like going outside to pick ya own switch.
luismartin757|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
luismartin757|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
ColorCated_Kita|odotkay|0.0|0.0|1.0|0.0|RT @odotkay: Just wanna know if Texas is gonna be District 8 or District 12 after this election. They might District 13 our asses.
peacelovespink|MannieMforever|-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
peacelovespink||-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
FerAmarante12|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
FerAmarante12|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
trimmgi|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
matslew|Slate|0.6808|0.0|0.682|0.318|Real time election projection by @Slate @Votecastr good decision and interesting journalistic experiment. https://t.co/YG88onihKi
matslew|slate|0.6808|0.0|0.682|0.318|Real time election projection by @Slate @Votecastr good decision and interesting journalistic experiment. https://t.co/YG88onihKi
DoctorBuxter|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
FireBox88|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
BettyBeene1|twitter|0.0|0.0|1.0|0.0|Election night at Huntsville Promenaders Square Dance Club. https://t.co/BPGZmYIDRb
DrBenz3|therealIRD|0.1832|0.121|0.725|0.154|RT @therealIRD: A brief break in my election obsession... to more normal obsession seeking justice in the #umc. https://t.co/t993SDFhSr
DrBenz3|twitter|0.1832|0.121|0.725|0.154|RT @therealIRD: A brief break in my election obsession... to more normal obsession seeking justice in the #umc. https://t.co/t993SDFhSr
nomadicdrift|bobfescoe|0.0|0.0|1.0|0.0|@bobfescoe we couldn't even figure out our own Brexit never mind the US election
hazucall|basket_mouth|0.0|0.0|1.0|0.0|@basket_mouth live on @TVCconnect. Speaking on US election https://t.co/SD18SAnHH0
hazucall|twitter|0.0|0.0|1.0|0.0|@basket_mouth live on @TVCconnect. Speaking on US election https://t.co/SD18SAnHH0
anya_fennec|theverge|0.3612|0.0|0.878|0.122|So there are a whole bunch of ways to stream the election news. Which ones do you guys like? https://t.co/AHJASRZy0l
trading24h|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
trading24h|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
SouthBeachSheed|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
SouthBeachSheed|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
DanielOzioma6|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
DanielOzioma6|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
knlaguerre|thetrudz|0.0|0.0|1.0|0.0|RT @thetrudz: 1) This is a long read. 2) This is personal. 3) Not debating a single word in it. 4) I think I am just about done discussing
Fanfan54T|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Fanfan54T|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
LibertyShaq|Cagsil|0.0382|0.0|0.943|0.057|@Cagsil then don't leave the house during any election or move to Cuba North Korea China or Qatar or something
DelawareFreedom|newsmax|0.0|0.0|1.0|0.0|RT @newsmax: Who are you voting for in this election? #MyVotes2016
adrijackson15|MissD4Trump|-0.4738|0.123|0.877|0.0|RT @MissD4Trump: This election will be decided by the people working 2 to 3 jobs.We need your vote! We need your evening vote! Ignore the T
RayLope20755050|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
QGS24|joe_fortkort5|0.1655|0.089|0.759|0.152|RT @joe_fortkort5: People love to talk about Hillary and Trump and how important this election is but forget the Warriors blew a 3-1 lead i
zoe_nor|latimes|0.0|0.0|1.0|0.0|"In Little Saigon, a possible generational divide at the polls https://t.co/PjvCdVmU0d"
carolrosenberg|MiamiHerald|0.0|0.0|1.0|0.0|@MiamiHerald newsroom fortifies for Election Night 2016. https://t.co/JkmkctQfQh
carolrosenberg|twitter|0.0|0.0|1.0|0.0|@MiamiHerald newsroom fortifies for Election Night 2016. https://t.co/JkmkctQfQh
bettyaberlin|Gabbienain|-0.6418|0.278|0.722|0.0|@Gabbienain this election has been so stressful for her she's going blonde.
ArlRooftop|WMALDC|0.4199|0.0|0.872|0.128|RT @WMALDC: We're ready to track the election state by state at Arlington Rooftop Bar and Grill! #ElectionNight #Election2016 https://t.co/
ArlRooftop|t|0.4199|0.0|0.872|0.128|RT @WMALDC: We're ready to track the election state by state at Arlington Rooftop Bar and Grill! #ElectionNight #Election2016 https://t.co/
viktoria_krolx|angusscottt|0.6369|0.0|0.822|0.178|RT @angusscottt: Canny wait for the American election to be over so we can focus on the real issues like if there's any hoose parties this
Margie71blue|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
awkksha|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
mlynne3|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
christhompson82|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
christhompson82|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
ToplessGoddess|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
ToplessGoddess|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
KristimoonAOA|instagram|-0.6597|0.293|0.707|0.0|"This has been such a draining and bizarre election season with that narcissistic, ego maniac, https://t.co/eD1J2bAvdV"
autobody65|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
stephanpippen|knbrmurph|-0.1531|0.06|0.94|0.0|RT @knbrmurph: Take a moment on Election Night to remember the Old School we all miss on TV: Big Tim Russert and the Magic Grease Board. #R
KevinJsAngels|deleasakathleen|0.0|0.0|1.0|0.0|@deleasakathleen this one? https://t.co/GErdcLVPcC
KevinJsAngels|m|0.0|0.0|1.0|0.0|@deleasakathleen this one? https://t.co/GErdcLVPcC
El4short|knbrmurph|-0.1531|0.06|0.94|0.0|RT @knbrmurph: Take a moment on Election Night to remember the Old School we all miss on TV: Big Tim Russert and the Magic Grease Board. #R
CorianderSleuth|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
CollectedN|latimes|0.0|0.0|1.0|0.0|Former President George W. Bush didn't vote for Donald Trump https://t.co/ZuKVSLGoH0
msdianesolomon|OPFergVal|-0.0571|0.131|0.71|0.159|RT @OPFergVal: So a large number of Trump supporters express their anger at @megynkelly and here she is to spoil election night on @foxnews
BigpapiHT|baratunde|0.0|0.0|1.0|0.0|RT @baratunde: So we are all watching Newsmax and Russia Today for the election results right?
DOOM2332|twitter|0.0|0.0|1.0|0.0|"Morrissey, on the Election- https://t.co/gXeYNo6i15"
BairdBev|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
distrumption|twitter|0.0|0.0|1.0|0.0|Thread #1  7:00pm Election Results and Discussion  #ElectionNight https://t.co/VlJ08cTt6F
viclyn529|WDFx2EU8|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
viclyn529|conservativeeagles|-0.7156|0.237|0.763|0.0|RT @WDFx2EU8: Breaking: Florida Election Worker Goes Public With Massive Voter Fraud Happening Right Now !!!!! https://t.co/m3jPrRGEXT
MexicanKeith|BeingKirst|0.0|0.0|1.0|0.0|@BeingKirst you should be more afraid of the election fo sho bro
amandalv845|twitter|0.0|0.0|1.0|0.0|This is what election night in the newsroom is all about #partylikeajournalist #workingtilmidnight https://t.co/QuA1YPdc8s
ScheeDawg|TheGoodGodAbove|-0.2263|0.087|0.913|0.0|"RT @TheGoodGodAbove: In 1996 Bob Dole fell off a stage not once, but twice.This election really could've used both candidates falling off"
kaylavelli|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
kaylavelli|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
bobbikitty|wolfieraps|0.7865|0.0|0.783|0.217|RT @wolfieraps: If trump wins the election today who wants to come back to Canada with me? LIKE this tweet so I know to buy you an airplane
Dougr6|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
Dougr6|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
AutumnAmadou|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
AutumnAmadou|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
venkyganesan|medium|0.7227|0.0|0.798|0.202|10 Things you will not read about in tomorrows papers but you should know regardless of who wins the election https://t.co/914cLjRffZ
ONLYTRUMP4USA|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
PeriodicaI|usatoday|0.197|0.0|0.861|0.139|Hillary Clinton calls voting for herself a 'most humbling feeling' - USA TODAY https://t.co/H70Ojke1Ob
gaboros|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
gaboros|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
The_Jodster_|natalieeecowann|-0.5719|0.227|0.773|0.0|RT @natalieeecowann: If you don't vote then you have no room to complain about how the election ends
GroverBeachBum|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
Christi0820|mike_pence|0.3818|0.0|0.894|0.106|"RT @mike_pence: The outcome of this historic election rests in your hands. If you stand for a stronger America, cast your vote for #TrumpPe"
lovelyVickyyy|_NisaJanaeee|0.5859|0.0|0.678|0.322|RT @_NisaJanaeee: If Trump win this election tonight https://t.co/vJJxm7efpZ
lovelyVickyyy|twitter|0.5859|0.0|0.678|0.322|RT @_NisaJanaeee: If Trump win this election tonight https://t.co/vJJxm7efpZ
sadmexicanchica|NathanZed|-0.25|0.215|0.601|0.184|RT @NathanZed: I remember back when this election was all fun and games like when we accused a candidate of being a serial murderer can we
krista_bach|SidneyCrosbyEgo|0.765|0.0|0.752|0.248|RT @SidneyCrosbyEgo: The best part about election day is that we get to watch McDavid and Crosby play before the world ends.
janettwokay|JoseAlmada_|0.3818|0.073|0.7|0.227|".@JoseAlmada_ Make sure to vote in every election, no matter how big or small it is, from here on out to eternity. Every vote matters. :-)"
rajuntexankajun|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
rajuntexankajun|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
Mr3lsewhere|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Mr3lsewhere|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
CollectedN|latimes|0.0|0.0|1.0|0.0|How this election has revealed workplace sexism is still an issue https://t.co/pGn0TMPnHa
WorldMktng|Queen_UK|0.5859|0.0|0.759|0.241|RT @Queen_UK: Very concerned that someone is going to win this election. #USElection
antfarmer|theaustralian|0.4927|0.0|0.834|0.166|Paul Kelly is very good here on Trump as a vandal and the decline of America ($) https://t.co/ydGRKhuvHc
MojoMelMM|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
MojoMelMM|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
pie_olaa|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
GermanT61734220|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
GermanT61734220|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
_Outerxspace|StephenKing|-0.34|0.103|0.897|0.0|"RT @StephenKing: The ugliest election in living memory is almost over, but the polls are still open. VOTE, PEOPLE. Do your job."
atticascott|funambulator|0.0|0.0|1.0|0.0|"RT @funambulator: Tune in to @WFPLNews 7-9pm for live election returns &amp; analysis with @atticascott, CW Julie Denton, @sean_southard &amp; @DSt"
sid4364|MannieMforever|-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
sid4364||-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
k8tlinbarajas|NathanZed|-0.25|0.215|0.601|0.184|RT @NathanZed: I remember back when this election was all fun and games like when we accused a candidate of being a serial murderer can we
scottt1984|steve68135|-0.5242|0.273|0.727|0.0|@steve68135 @DebAlwaystrump @stmpinfortrump A bunch of lies! Obama rigging the election!
Inked_Banana|politico|0.0|0.0|1.0|0.0|"RT @politico: #BREAKING: Results of the U.S. elections are beginning to flow in, starting with returns from Indiana and Kentucky https://t."
Inked_Banana||0.0|0.0|1.0|0.0|"RT @politico: #BREAKING: Results of the U.S. elections are beginning to flow in, starting with returns from Indiana and Kentucky https://t."
piimavaras|Night_0f_Fire|-0.4574|0.286|0.549|0.165|Mass shooter #SamHyde is active again and killing voters! https://t.co/OHzMIrWktU @Night_0f_Fire
piimavaras|rt|-0.4574|0.286|0.549|0.165|Mass shooter #SamHyde is active again and killing voters! https://t.co/OHzMIrWktU @Night_0f_Fire
MacDHistory|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: The latest updates on the House races https://t.co/Q1iwJbI6El https://t.co/SvkRA88ctf
MacDHistory|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: The latest updates on the House races https://t.co/Q1iwJbI6El https://t.co/SvkRA88ctf
hopi2lotus|900amWURD|0.3595|0.0|0.906|0.094|RT @900amWURD: We're live at @EnonTab for the rest of Election Night! Join us at 2800 W. Cheltenham Ave. to watch results come in. https://
hopi2lotus||0.3595|0.0|0.906|0.094|RT @900amWURD: We're live at @EnonTab for the rest of Election Night! Join us at 2800 W. Cheltenham Ave. to watch results come in. https://
ShebaJo|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
ShebaJo|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
amityville315x|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
gascasf|Twitter|0.0|0.0|1.0|0.0|Election coverage on Twitter @Twitter https://t.co/OvHVLY9jdn
gascasf|twitter|0.0|0.0|1.0|0.0|Election coverage on Twitter @Twitter https://t.co/OvHVLY9jdn
MargHartmann|vox|0.357|0.0|0.84|0.16|As if I werent jealous enough that my polling place doesnt do I voted stickers https://t.co/Kf8XoPXTpG
Joanne1009|CNN|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
Joanne1009|twitter|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
TheMowll|jerome_corsi|-0.5859|0.153|0.847|0.0|RT @jerome_corsi: TRUMP NEEDS ALL POSSIBLE VOTERS IN PA - voter fraud being reported EVENING HOURS WILL DECIDE ELECTION - get all Trump vot
Magitroopa|CBSThisMorning|0.0|0.0|1.0|0.0|RT @CBSThisMorning: Oh how this map will change. How Election night begins... #CBSElection  https://t.co/SraM591OGV
Magitroopa|twitter|0.0|0.0|1.0|0.0|RT @CBSThisMorning: Oh how this map will change. How Election night begins... #CBSElection  https://t.co/SraM591OGV
bookbeaut|twitter|-0.5983|0.251|0.659|0.091|"Combating election anxiety by replying to emails from this experiment tonight! Come, join, tell me the worst time y https://t.co/I5ra1X5dZI"
flicofthetongue|BuzzFeedNews|0.3595|0.0|0.884|0.116|RT @BuzzFeedNews: The  time  has  come! Join BuzzFeed News LIVE on Twitter as we get through #ElectionNight results together  https://
flicofthetongue||0.3595|0.0|0.884|0.116|RT @BuzzFeedNews: The  time  has  come! Join BuzzFeed News LIVE on Twitter as we get through #ElectionNight results together  https://
RichSuchet|iandstone|0.0|0.0|1.0|0.0|@iandstone I just had a look to see what's really happening out there. It turns out the US election is a sideshow: https://t.co/O1emNtLc4L
RichSuchet|twitter|0.0|0.0|1.0|0.0|@iandstone I just had a look to see what's really happening out there. It turns out the US election is a sideshow: https://t.co/O1emNtLc4L
MarieCamalier|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
MarieCamalier|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
jjnado|MikeDrucker|0.0|0.0|1.0|0.0|RT @MikeDrucker: Yo can we have a big smash bros tournament on your screens after the election https://t.co/Zda4wZIh88
jjnado|twitter|0.0|0.0|1.0|0.0|RT @MikeDrucker: Yo can we have a big smash bros tournament on your screens after the election https://t.co/Zda4wZIh88
ChiefKota_TYB|Yike4Tyke|0.4215|0.0|0.859|0.141|"@Yike4Tyke she also has 0.3% of the popular vote, the same percentage she had in the 2012 election"
MelodyTruong|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
MelodyTruong|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
elaine_wildes|asdomke|-0.6249|0.282|0.718|0.0|RT @asdomke: Polls disappear showing major Hillary collapse among likely voters on election day... https://t.co/zI3JeNYMCO
elaine_wildes|linkis|-0.6249|0.282|0.718|0.0|RT @asdomke: Polls disappear showing major Hillary collapse among likely voters on election day... https://t.co/zI3JeNYMCO
JamesTricePPP|IamJasonSole|0.0|0.0|1.0|0.0|"RT @IamJasonSole: Waiting a long time to vote in a presidential election! I did it for the 51,000 disenfranchised.#RestoretheVoteMN https:"
sandimac|vermontgmg|0.0|0.0|1.0|0.0|"RT @vermontgmg: As the first major set of polls close, here's what the data nerds will be watching as the results come in: https://t.co/TI0"
sandimac|t|0.0|0.0|1.0|0.0|"RT @vermontgmg: As the first major set of polls close, here's what the data nerds will be watching as the results come in: https://t.co/TI0"
AGuercy|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
AGuercy|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
kriketUSA|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
kriketUSA|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
Ayooo_Serenity|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
Ayooo_Serenity|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
Raveneyes|untappd!|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/u2KvtVXd7d #voteforbeer
Raveneyes|untappd|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/u2KvtVXd7d #voteforbeer
abs_tellthetale|dorseyshaw|0.0|0.0|1.0|0.0|RT @dorseyshaw: I think Chris Matthews just said Tip O'Neill and JFK went to a porn theater on Election Night back in the day https://t.co/
abs_tellthetale|t|0.0|0.0|1.0|0.0|RT @dorseyshaw: I think Chris Matthews just said Tip O'Neill and JFK went to a porn theater on Election Night back in the day https://t.co/
skohayes|DrDigiPol|0.4574|0.0|0.813|0.187|RT @DrDigiPol: Trump opts to have his election funeral... err... party at a unionized hotel!#ElectionNight
flmabon|instagram|0.5719|0.0|0.654|0.346|Yup this just happened.  Happy Election 2016 https://t.co/t8mhways3H
vavoida|AnnLe__|0.25|0.0|0.667|0.333|@AnnLe__ gonna be alright https://t.co/8ZhDXM3rzv
vavoida|ianwelsh|0.25|0.0|0.667|0.333|@AnnLe__ gonna be alright https://t.co/8ZhDXM3rzv
_FaisalSayed|Telegraph|-0.6486|0.223|0.777|0.0|RT @Telegraph: #ElectionNight One person is reportedly dead after a shooting in California near a polling station https://t.co/CJCBsKKKNE
_FaisalSayed|telegraph|-0.6486|0.223|0.777|0.0|RT @Telegraph: #ElectionNight One person is reportedly dead after a shooting in California near a polling station https://t.co/CJCBsKKKNE
pendekarsilat11|Myrmecos|0.6124|0.11|0.596|0.294|RT @Myrmecos: We interrupt your election to bring you a yellow butterfly of peace and hope. https://t.co/RVbcdKeYsa
pendekarsilat11|twitter|0.6124|0.11|0.596|0.294|RT @Myrmecos: We interrupt your election to bring you a yellow butterfly of peace and hope. https://t.co/RVbcdKeYsa
HashtagGrateful|kstlz|0.4588|0.0|0.88|0.12|RT @kstlz: 2day Im grateful for my ID which allowed me 2 vote 2day &amp; buy election recovery booze after #grateful #ThxObama #literallytho #u
simonvandore|insightSBS|0.0|0.0|1.0|0.0|RT @insightSBS: Follow the votes as they roll in from today's momentous US Presidential Election: https://t.co/ralz3v4M0E @SBSNews https://
simonvandore|sbs|0.0|0.0|1.0|0.0|RT @insightSBS: Follow the votes as they roll in from today's momentous US Presidential Election: https://t.co/ralz3v4M0E @SBSNews https://
keen_kyungsoo|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
keen_kyungsoo|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
bestpartyleon|mashable|0.0|0.0|1.0|0.0|America gets lit: The Lite Brite guide to election results https://t.co/TwBBkJJQOj
MattyDHarris784|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
MattyDHarris784|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
JuliaInLights|MattBellassai|-0.0258|0.131|0.742|0.127|"RT @MattBellassai: hey @realDonaldTrump just wanna say that despite everything that's happened this election, you're still awful and i hope"
fluffynutters|Jonbuckhouse|0.6239|0.0|0.843|0.157|RT @Jonbuckhouse: The Polls are starting to close all over the US! Who do you think will win the election?  #ElectionNight #electionday #iV
JackJrl935|mike_pence|0.0|0.0|1.0|0.0|"RT @mike_pence: This Election Day, America is standing at the crossroads of history. RT this if you're voting for @realDonaldTrump. Togethe"
angelacdumlao|fakedansavage|-0.2579|0.165|0.733|0.102|RT @fakedansavage: I'm retweeting a Republican without sarcasm or snark - this election is insane. https://t.co/mvaoZO0elr
angelacdumlao|twitter|-0.2579|0.165|0.733|0.102|RT @fakedansavage: I'm retweeting a Republican without sarcasm or snark - this election is insane. https://t.co/mvaoZO0elr
hopelmez16|dougsmith1946|0.0|0.0|1.0|0.0|RT @dougsmith1946: @nationdivided @janiehburton  @FBI @FBIWFO  @NewYorkFBI  That's why officials stuffed ballot boxes for Hillary https://t
hopelmez16||0.0|0.0|1.0|0.0|RT @dougsmith1946: @nationdivided @janiehburton  @FBI @FBIWFO  @NewYorkFBI  That's why officials stuffed ballot boxes for Hillary https://t
castraley|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
aacoek|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
aacoek|t|0.0|0.0|1.0|0.0|RT @wikileaks: Assange statement: What are the reasons behind WikiLeaks exposures of the DNC and the Clinton campaign? https://t.co/Q6KEChq
usa67us|EdBaker3000|0.2263|0.0|0.863|0.137|RT @EdBaker3000: Officials: PA Voting Machines Incorrectly Registered Straight Republican Votes - Breitbart https://t.co/FVcPeTI6FE
usa67us|breitbart|0.2263|0.0|0.863|0.137|RT @EdBaker3000: Officials: PA Voting Machines Incorrectly Registered Straight Republican Votes - Breitbart https://t.co/FVcPeTI6FE
rosegoggles|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
rosegoggles|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
jwead4570|pmicc33|0.555|0.106|0.636|0.258|"RT @pmicc33: Soros strikes again!Keep it up losers,you'll invalidate the whole election.Trump supporters will only accept a Trump win!#M"
cheryl_hardt|mw_bizwomen|0.4404|0.0|0.861|0.139|RT @mw_bizwomen: Need a break from election coverage? Read how @CREW_Network is building a better pipeline in commercial real estate https:
joelsblankspace|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
joelsblankspace|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
blujaydavid|LaurenJauregui|0.4795|0.0|0.881|0.119|RT @LaurenJauregui: I'm so excited that I was able to exercise my vote as a Cuban American Woman for the first time in this particular elec
imranmeyan|GAVlNREACTS|0.6249|0.0|0.661|0.339|RT @GAVlNREACTS: A great way to start Election Day https://t.co/yr6QAP3orF
imranmeyan|twitter|0.6249|0.0|0.661|0.339|RT @GAVlNREACTS: A great way to start Election Day https://t.co/yr6QAP3orF
JasonAmessenger|twitter|0.0|0.0|1.0|0.0|Obligatory Election Night tweet https://t.co/43QwBDvDfX
FreshDialogues|nytimes|0.5859|0.0|0.725|0.275|RT @nytimes: When will we know when we have a winner? https://t.co/58YOEs664i
FreshDialogues|nytimes|0.5859|0.0|0.725|0.275|RT @nytimes: When will we know when we have a winner? https://t.co/58YOEs664i
EidojTrump|TheLastRefuge2|0.0|0.0|1.0|0.0|RT @TheLastRefuge2: Thread #1  7:00pm Election Results and Discussion https://t.co/dvp9W1yfpJ https://t.co/1kuDOKqQA4
EidojTrump|theconservativetreehouse|0.0|0.0|1.0|0.0|RT @TheLastRefuge2: Thread #1  7:00pm Election Results and Discussion https://t.co/dvp9W1yfpJ https://t.co/1kuDOKqQA4
JaimeHdezAmin|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
JaimeHdezAmin|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
TerryLeeUSA|politico|0.0|0.0|1.0|0.0|Live Map is Up https://t.co/wtRieFM0yl
FightingTories|ABCaustralia|-0.7845|0.317|0.683|0.0|Bloody childish and trash coverage as the @ABCaustralia @abcnews24 waste taxpayer dollars on the US election. The Guthrie factor #ABCTRASHED
MHB1070|ForTrump|0.3182|0.0|0.909|0.091|RT @ForTrump: Please get out and vote. Do not listen 2exit polls. This is the election that will decide our country's future.  Let's #MAGA
JessieJessie08|JMick1734|0.0|0.0|1.0|0.0|RT @JMick1734: This election reminds me of dan scott vs karen rowe when they ran for mayor of tree hill
lauren_detrich|Max_Shores20|0.0|0.0|1.0|0.0|RT @Max_Shores20: #MannequinChallenge Election Day Purge theme! https://t.co/C6Oxgr0xPi
lauren_detrich|twitter|0.0|0.0|1.0|0.0|RT @Max_Shores20: #MannequinChallenge Election Day Purge theme! https://t.co/C6Oxgr0xPi
peterbilt00|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you VOTED TO DRAIN THE SWAMP! #MAGA #ElectionDay #Election https://t.co/TkUPGBNYkg
peterbilt00|twitter|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you VOTED TO DRAIN THE SWAMP! #MAGA #ElectionDay #Election https://t.co/TkUPGBNYkg
AlisonVerhoeven|twitter|0.0|0.0|1.0|0.0|All dressed up in Washington for election night #USTour https://t.co/ckeCWt0OQs
NWONightmare|TrumpWinner_16|-0.6884|0.226|0.774|0.0|RT @TrumpWinner_16: Florida Election Worker Went Public With Massive Voter Fraud GOING DOWN RIGHT NOW!!! https://t.co/m8z2QeXlaR https://t.
NWONightmare|everynewshere|-0.6884|0.226|0.774|0.0|RT @TrumpWinner_16: Florida Election Worker Went Public With Massive Voter Fraud GOING DOWN RIGHT NOW!!! https://t.co/m8z2QeXlaR https://t.
FilipDobi|SebGorka|0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
FilipDobi||0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
JDE6321|realDonaldTrump|0.0|0.0|1.0|0.0|"RT @realDonaldTrump: Before my FINAL campaign speech, I will get a list of Election Day Donors! Donate NOW! https://t.co/iZjo4q2gYA https:/"
JDE6321|secure|0.0|0.0|1.0|0.0|"RT @realDonaldTrump: Before my FINAL campaign speech, I will get a list of Election Day Donors! Donate NOW! https://t.co/iZjo4q2gYA https:/"
TiffanyRothe|youtube|0.0|0.0|1.0|0.0|Don't be the one with excuses. This election is bigger than the candidates. https://t.co/FZF06ODW3l
breedloveme|heywtfabi|-0.5994|0.495|0.505|0.0|@heywtfabi too anxious abt election results :(
GeorgeJB1990|twitter|0.8475|0.0|0.566|0.434|"Tonight's election is a lot like 'Alien vs Predator', 'Whoever wins, we loose'! Ha! #Truth4751 https://t.co/VaqgmSe79q"
KarinMStone|drsteuss|0.6369|0.0|0.802|0.198|RT @drsteuss: The merch is ready to go at the DFL election party. More election coverage coming up on @kare11 at 6. https://t.co/lWBY0KVky1
KarinMStone|twitter|0.6369|0.0|0.802|0.198|RT @drsteuss: The merch is ready to go at the DFL election party. More election coverage coming up on @kare11 at 6. https://t.co/lWBY0KVky1
kinshasaweb|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
kinshasaweb|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
HadleyKiefer|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
HadleyKiefer|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
NECN|necn|0.0|0.0|1.0|0.0|WATCH LIVE: necn's election night coverage. https://t.co/TjMPutYNa0
caseyyy_h|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
caseyyy_h|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
whynotmeplease|SavidgeReads|0.5994|0.0|0.824|0.176|"RT @SavidgeReads: Dear Santa, as an early Christmas present please let me wake up to the election of the first female president of the USA."
kid_twist|_alastair|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
kid_twist|t|0.624|0.0|0.796|0.204|RT @_alastair: The @GuardianUS interactive team has a really amazing map display for tonight's results. Take a look: https://t.co/hFTmGzGAr
alexn_leigh|dril|0.0|0.0|1.0|0.0|RT @dril: if you ask me this election could end about 100 different ways:1) trump gets 0% of the vote2) trump gets 1% of the vote3) trum
threestangtyry|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
_tyler_tyler|JohnKingCNN|0.4019|0.0|0.847|0.153|I wish to one day thrive in my life the way @JohnKingCNN thrives at the Election SmartBoard.
OakvilleDad|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
OakvilleDad|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
_lowkeymaya|maitlynxo|-0.5319|0.135|0.865|0.0|RT @maitlynxo: If you are 18+ and didn't vote I don't wanna hear NA COMPLAINTS about the election because you didn't do your part.
JoshCovitt|ucbtla|0.0|0.0|1.0|0.0|RT @ucbtla: $5 #ElectionDay shows at @ucbsunset https://t.co/OKj0Ren3CY7pm Election Scenes 8:30pm Election Results Live 10:30pm Outsi
JoshCovitt|t|0.0|0.0|1.0|0.0|RT @ucbtla: $5 #ElectionDay shows at @ucbsunset https://t.co/OKj0Ren3CY7pm Election Scenes 8:30pm Election Results Live 10:30pm Outsi
ibickis|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
lisamakela2|WordSmithGuy|0.0|0.0|1.0|0.0|RT @WordSmithGuy: Florida Panhandle &amp; Michigan: You have 1 hour &amp; 15 minutes to make history. This entire election may be decided by you gu
shaveblog|nytimes!https//t.co/dEpEujj534|0.0|0.0|1.0|0.0|"Heckuva job, @nytimes!https://t.co/dEpEujj534"
shaveblog|nytimes|0.0|0.0|1.0|0.0|"Heckuva job, @nytimes!https://t.co/dEpEujj534"
jcmenacho93|nytopinion|0.0|0.0|1.0|0.0|RT @nytopinion: The too long 2016 campaign ends when you vote in today's election. And then: we hold our breath. https://t.co/TKzCHO2BLk ht
jcmenacho93|nytimes|0.0|0.0|1.0|0.0|RT @nytopinion: The too long 2016 campaign ends when you vote in today's election. And then: we hold our breath. https://t.co/TKzCHO2BLk ht
centroarsnatur1|centroarsnatura|0.0|0.0|1.0|0.0|"""How the Pro-Trump Media Covered Election Day"" by JOHN HERRMAN and SAPNA MAHESHWARI via NYT  https://t.co/Khhg46LV6E"
ShawnPoss|SebGorka|0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
ShawnPoss||0.8779|0.0|0.558|0.442|"RT @SebGorka: Good sign:Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' https://t."
JasmineAyadova|ddlovato|0.1027|0.101|0.734|0.165|RT @ddlovato: I apologize for the joke I made earlier.. seemed to offend some people. Just making light of the election 
Stevepppppppp|cnbc|0.0|0.0|1.0|0.0|"Showdown in the Buckeye State: 'As Ohio goes, so goes the nation' https://t.co/gOtap2L6AI #Election2016"
9NEWS|9news|0.2023|0.135|0.676|0.189|Stuck in a line to vote? Here some entertainment while you wait: https://t.co/PQcmFhmWv7
theledger|madisonfantozzi|0.4019|0.0|0.876|0.124|RT @madisonfantozzi: My first #electiondaypizza ever. Yes I've worked in newsrooms for 4+ years... this election I've been #blessed https:/
theledger||0.4019|0.0|0.876|0.124|RT @madisonfantozzi: My first #electiondaypizza ever. Yes I've worked in newsrooms for 4+ years... this election I've been #blessed https:/
FYC_Crow|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
FYC_Crow|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
UCentralMedia|facebook|0.0|0.0|1.0|0.0|UCentral Election 2016 https://t.co/5edphDFLJe
naomibeast_|WORLDSTAR|0.5859|0.0|0.678|0.322|RT @WORLDSTAR: Who will win the 2016 presidential election? 
shrynyk|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
NickDawybida|ConanOBrien|0.8271|0.0|0.7|0.3|RT @ConanOBrien: Congratulations to the winner of the 2016 presidential election.  Youll be receiving the cleaning bill for Americas pant
ashleyavila_|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
margimcclelland|TheLastRefuge2|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
margimcclelland|twitter|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
1isten_up|dcexaminer|0.0|0.0|1.0|0.0|RT @dcexaminer: The first polls in Florida are about to close. Full state closings and our live electoral map: https://t.co/Iz2vhOwGcW #Ele
1isten_up|washingtonexaminer|0.0|0.0|1.0|0.0|RT @dcexaminer: The first polls in Florida are about to close. Full state closings and our live electoral map: https://t.co/Iz2vhOwGcW #Ele
welcome_2KBToys|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
welcome_2KBToys|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
chrishuff_sf|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
bblancoynot|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
profmusgrave|CNN|0.0|0.0|1.0|0.0|"Our election night plan: @CNN , alcohol, and Middle Eastern cuisine."
halogalopagos|SarahCAndersen|-0.1531|0.086|0.914|0.0|RT @SarahCAndersen: Need to finish tomorrow's comic but the election is messing with my nerves just a LITTLE https://t.co/XjkCcpqXsV
halogalopagos|twitter|-0.1531|0.086|0.914|0.0|RT @SarahCAndersen: Need to finish tomorrow's comic but the election is messing with my nerves just a LITTLE https://t.co/XjkCcpqXsV
PatriotCzar|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
HatokTalk|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
efm6660|instagram|0.0|0.0|1.0|0.0|"Election Night 2016. TV on, pumpkin carved. #election2016 #electionnight https://t.co/IF03pDGZuD"
CollectedN|cnn|0.0|0.0|1.0|0.0|"Control of Senate, House up for grabs https://t.co/U1jcF8nCXQ"
GerikaTurner|cuddlereedus|0.6654|0.0|0.611|0.389|RT @cuddlereedus: vote! who should win the election??
tvheidihatch|twitter|0.4404|0.0|0.854|0.146|Good plan. I remember my 1st presidential election. The Presidential race had been called before I cast my ballot.  https://t.co/DfFk1bI9jc
upflund|naonaophoto|0.5538|0.0|0.826|0.174|RT @naonaophoto: It's interesting to see such variety perspectives towards the US election via this event tonight!!! #usewlund
stuart_goldman|twitter|0.0|0.0|1.0|0.0|Every Friday night is an election night for high school sports at a newspaper. https://t.co/8tLnn9zcV0
LeslieWix|CBSNews|0.2716|0.0|0.909|0.091|RT @CBSNews: First exit poll of Election 2016 shows that the most important issue to North Carolina is the economy #Election2016 https://t.
LeslieWix||0.2716|0.0|0.909|0.091|RT @CBSNews: First exit poll of Election 2016 shows that the most important issue to North Carolina is the economy #Election2016 https://t.
johnnykats|FiveThirtyEight|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
johnnykats|t|0.6908|0.087|0.655|0.258|"RT @FiveThirtyEight: If Clinton wins Florida, her probability of winning the Electoral College would shoot up to 93% from 71%. https://t.co"
MicahKool|TheRock|0.0|0.0|1.0|0.0|"This has to be the first election ever where more people ask you ""who'd you write in?"" Instead of ""who'd you vote for?"" My answer: @TheRock"
katelynd_hill87|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
joeldoesnothing|Angryish|0.8008|0.043|0.699|0.259|"@Angryish I never want to hear about this election again. Ever. Let's talk about fun things. Cats, dogs, video games, how great Joel is..."
Meganwiley204|mitchellvii|0.5267|0.0|0.848|0.152|"RT @mitchellvii: Democracy Institute, ONLY pollster to correctly guess Brexit, has Trump winning by 5.  Same as my prediction:  https://t.c"
Meganwiley204||0.5267|0.0|0.848|0.152|"RT @mitchellvii: Democracy Institute, ONLY pollster to correctly guess Brexit, has Trump winning by 5.  Same as my prediction:  https://t.c"
rebekka_jf|fromrosesxo|-0.067|0.088|0.836|0.077|RT @fromrosesxo: I know I'm not alone when I say I've got anxious Brexit type feelings again about the result of the election.
KaitlynHalfPint|BradyHaran|0.0|0.094|0.812|0.094|"RT @BradyHaran: No joke, hardest thing about following US election coverage is remembering that red means Republican &amp; blue means Democrat."
liyuanwei|qz|0.0|0.0|1.0|0.0|RT @qz: From Nina Simone to Beyonce: The Quartz playlist of songs by women who rule https://t.co/34y9D4BdxT
liyuanwei|qz|0.0|0.0|1.0|0.0|RT @qz: From Nina Simone to Beyonce: The Quartz playlist of songs by women who rule https://t.co/34y9D4BdxT
JohnTuckah|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
deachterdeur|vocnederland|0.0|0.0|1.0|0.0|RT @vocnederland: Live Cannabis Legalization Coverage &amp; Results: Election 2016 | Leafly https://t.co/tqWv3lPO7A #cannabis #leafly via @Leaf
deachterdeur|leafly|0.0|0.0|1.0|0.0|RT @vocnederland: Live Cannabis Legalization Coverage &amp; Results: Election 2016 | Leafly https://t.co/tqWv3lPO7A #cannabis #leafly via @Leaf
efairhurst|digitaltrends|0.0|0.0|1.0|0.0|"How to track the 2016 election results with every map, graph, and poll online https://t.co/WoLjKOwTw0"
MadHermit|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
MadHermit|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
vrai777|bloomberg|0.0|0.0|1.0|0.0|#BloombergTV  We're live-blogging #ElectionNight results. Follow along here https://t.co/OV4nr2UhZY https://t.co/QGTVBjImiG
Smedley_Butler|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Election Results #ElectionDay https://t.co/fBR9hVgWHg
Smedley_Butler|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Election Results #ElectionDay https://t.co/fBR9hVgWHg
CndnDwnSouth|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
TimerUsa|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
TimerUsa|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
MichaelBarger1|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
MichaelBarger1|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
Dadspar|twitter|0.5106|0.0|0.82|0.18|"Bill's earnest tweets are the only thing keeping me sane in this zany election, folks. https://t.co/ZEbt2FT6T5"
TonyBeavers1|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
Cediwaa|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
Cediwaa|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
SoCalPhillie|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
clrih9|Millican21|0.0|0.0|1.0|0.0|RT @Millican21: Getting my election coverage from @SamSeder and @_michaelbrooks on the @majorityfm YouTube channel.
boyzer23|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
boyzer23|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
ash00200|ABC7Chicago|0.25|0.0|0.917|0.083|RT @ABC7Chicago: Chance the Rapper leads hundreds of young voters to long early voting lines downtown so they can cast their ballots: https
JohnZorabedian|CraigSilverman|-0.4767|0.147|0.853|0.0|RT @CraigSilverman: New debunks: Soros-connected voting machines are NOT being used today Beware of a fake CNN Politics account http
Aupps|untappd!|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/Q6uKZv1Bzt #voteforbeer
Aupps|untappd|0.0|0.0|1.0|0.0|I just earned the 'Election Day (2016)' badge on @untappd! https://t.co/Q6uKZv1Bzt #voteforbeer
MonroesMindset|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
OMHSmedia|nprpolitics|0.0|0.0|1.0|0.0|"RT @nprpolitics: For full coverage and analysis, follow our live blog. https://t.co/0WfRXoXnye #ElectionDay #Election2016 https://t.co/Rcqe"
OMHSmedia|npr|0.0|0.0|1.0|0.0|"RT @nprpolitics: For full coverage and analysis, follow our live blog. https://t.co/0WfRXoXnye #ElectionDay #Election2016 https://t.co/Rcqe"
FLady37m|hrtablaze|0.9207|0.0|0.645|0.355|RT @hrtablaze: My Bernie Sanders loving nephew who has been messing with me all election just told me he voted TRUMP !!! WOOT WOOT ! #elect
ulilgypsy|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
ulilgypsy|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
MuzikMan1977|MuzikMan1977|0.0|0.0|1.0|0.0|"RT @MuzikMan1977: This is my ""2016 Election Command Center"" #vote #election2016 #Technology #cyber #polls #bigdata #exitpolls #CNN #MSNBC #"
CarolynGambon|MannieMforever|-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
CarolynGambon||-0.8979|0.459|0.541|0.0|"RT @MannieMforever: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
motherthot|carwash54|0.7085|0.0|0.734|0.266|"RT @carwash54: Me @ the beginning of the election: Ain't no way America letting a cheeto become president. lol what a joke Me November 7,"
wanthillaryout|twitter|0.0|0.0|1.0|0.0|realDenaldTrump: RT Harringtonkent: Here's the most insightful (and funny) pundit this election cycle https://t.co/qqs6qrUX3K
ktnote|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
ktnote|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
jjbaker333|CBCAlerts|-0.8481|0.326|0.674|0.0|"RT @CBCAlerts: One dead in shooting in California, three injured near polling station. No indication so far that it is election-related: re"
Bolopion|samueloakford|0.9344|0.0|0.497|0.503|RT @samueloakford: A bit of non-election news: deeply honored and grateful to have been awarded the @unfoundation's top prize for humanitar
raphaellaN|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
raphaellaN|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Basi20|Phil_Lewis_|-0.296|0.136|0.864|0.0|RT @Phil_Lewis_: These black women also deserve a visit to their graves on #ElectionDay https://t.co/8s4oXZTCvQ https://t.co/4opePa8GKg
Basi20|huffingtonpost|-0.296|0.136|0.864|0.0|RT @Phil_Lewis_: These black women also deserve a visit to their graves on #ElectionDay https://t.co/8s4oXZTCvQ https://t.co/4opePa8GKg
RichardDBK|RichardDBK|-0.2732|0.091|0.864|0.045|"@RichardDBK No matter what you think of Hillary, that should at least give you pause to think about how historic this election is."
firetomfriedman|politico|-0.4767|0.147|0.853|0.0|Clinton couldn't even wait for polls to close to rub our noses in how fake the election was. https://t.co/ykWC3xmx56
AnyonebutConnor|theJeremyVine|0.0|0.0|1.0|0.0|You know it's an election night when @theJeremyVine gets his multicoloured graphics out.
reneegoldsbery|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
frankzulla|DiamondGirl127|0.2732|0.077|0.807|0.116|"RT @DiamondGirl127: Voting monitor: Weren't you here earlier?Me: Uh no. Trust me lady, the last thing I'm trying to do is vote twice in th"
jefferymonaghan|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
steve2noriko|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
steve2noriko||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
esquire|ESQPolitics|0.6369|0.0|0.606|0.394|RT @ESQPolitics: They're ready to party in Philadelphia https://t.co/j4XQCQ7pTz https://t.co/EPyxA2ODgD
esquire|esquire|0.6369|0.0|0.606|0.394|RT @ESQPolitics: They're ready to party in Philadelphia https://t.co/j4XQCQ7pTz https://t.co/EPyxA2ODgD
DrKevGuitar|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
Chloe2229|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
heeyitsSJ|hannahjewcy|0.0|0.0|1.0|0.0|Thinking of @hannahjewcy and all others in the USA who have been so triggered by this election
z4mp1|blog|0.5106|0.0|0.87|0.13|Sling: Hey_Landon We still have the channels here on Sling TV. You can try us out by signing up for tonight's free https://t.co/LtBv3L1lfd
SithAlkline|champagnepapi|0.5719|0.0|0.791|0.209|RT @champagnepapi: If Donald trump wins the election I'll PayPal everyone that rted this $1
mckennaa_dugan|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
mckennaa_dugan|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
cnbintucson|JJohnsonLaw|-0.1531|0.18|0.67|0.149|@JJohnsonLaw @azmoderate I hope that guy ends up with a felony conviction and can't vote next election.
jaackiiee_o|instagram|0.0|0.0|1.0|0.0|"Election Night ritual since I was 8 yrs old: dad, me, nat'l news, KET, local radio updates, and https://t.co/9WMz6Y8J0J"
AAbramshe|MrMikeCalta|0.8165|0.0|0.616|0.384|So awesome to hear @MrMikeCalta  and @DrewOnTheRadio!  Thank you for the election coverage! #Election2016
efairhurst|latimes|0.0|0.0|1.0|0.0|Election day 2016 live updates: Early results are now coming in https://t.co/LAo87iih0b
lukestrat14|ESPNStatsInfo|0.34|0.0|0.906|0.094|RT @ESPNStatsInfo: Connor McDavid &amp; Sidney Crosby meet for 1st timeMario Lemieux &amp; Wayne Gretzky played vs each other for 1st time on Ele
RHS_APecon|WSJecon|0.3182|0.104|0.736|0.16|"RT @WSJecon: If Donald Trump wins, stock markets will likely fall and uncertainty will rise, Greg Ip writes https://t.co/IeKbqTQOGv "
RHS_APecon|blogs|0.3182|0.104|0.736|0.16|"RT @WSJecon: If Donald Trump wins, stock markets will likely fall and uncertainty will rise, Greg Ip writes https://t.co/IeKbqTQOGv "
radiojosie|FireballWhisky|0.0|0.0|1.0|0.0|Election Day coverage... @FireballWhisky or @BulleitUSA #rye #whiskey 
CassellCaptain|twitter|0.4404|0.0|0.775|0.225| if you need something to brighten your Election Day #Hokies https://t.co/KCADwtpoKw
ariiimichelle|kaiiclayy|-0.3605|0.177|0.699|0.124|"RT @kaiiclayy: this election has brought nothing but negativity and hate towards one another, we need a president who's going to bring noth"
panarmstrong|midcitymessenger|0.0|0.0|1.0|0.0|"Meanwhile in New Orleans, it is just another Tuesday election (because we have a lot of elections). #NOLA #GeauxVote https://t.co/V7w0VjC3RX"
wolvesmasks|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
wolvesmasks|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
WolfsonLiterary|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
WolfsonLiterary|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
SandieHelm|pmicc33|-0.7035|0.273|0.654|0.072|"RT @pmicc33: If we haven't learned anything in this election,1 thing is definite, the Democrats are a bunch of cheaters who cannot win fair"
__cassidyharris|bholtvluwer|0.8881|0.0|0.572|0.428|RT @bholtvluwer: Election Day fun with @GoNoodle ! Thank you #BlazerFresh for an awesome song!  #votevotevote  #cwcline https://t.co/Em3O
__cassidyharris|t|0.8881|0.0|0.572|0.428|RT @bholtvluwer: Election Day fun with @GoNoodle ! Thank you #BlazerFresh for an awesome song!  #votevotevote  #cwcline https://t.co/Em3O
JustMe725|ozarkadian|0.0|0.0|1.0|0.0|"RT @ozarkadian: #NoSleepTilPOTUS  OMG I swore I wouldn't follow the election results, but here I am -- watching. https://t.co/gR4CFyHbMY"
JustMe725|twitter|0.0|0.0|1.0|0.0|"RT @ozarkadian: #NoSleepTilPOTUS  OMG I swore I wouldn't follow the election results, but here I am -- watching. https://t.co/gR4CFyHbMY"
ThomasAHester2|spkhp|0.296|0.0|0.872|0.128|"RT @spkhp: Me: Who are you voting for in the election?1st grader: My momMe: Yeah, same"
dianuuhh|REALBrianStreng|0.7096|0.0|0.789|0.211|RT @REALBrianStreng: Joke is on Hillary if she wins the election because that means she has to sit at the desk Monica was under
USA_with_Trump|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
notsurewhere|layingbackeatin|-0.5106|0.268|0.732|0.0|RT @layingbackeatin: #ElectionDay I am actually physically sick of this election.
Grant_Robinson1|ZachAJacobson|0.0|0.0|1.0|0.0|RT @ZachAJacobson: Election Day reminder not to let political stance/indifferences:1. Define you.2. Get in the way of any personal relati
bbttttttt|GoAngelo|0.0|0.0|1.0|0.0|"RT @GoAngelo: Election Night 2012Actual ResultsObama: 65,915,795Romney: 60,933,504 https://t.co/dtD8WwpAd6"
bbttttttt|twitter|0.0|0.0|1.0|0.0|"RT @GoAngelo: Election Night 2012Actual ResultsObama: 65,915,795Romney: 60,933,504 https://t.co/dtD8WwpAd6"
scottpadair|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
AmeliaO28929509|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: Kai sporting the #MAGA hat. She has only asked 300 times today if she could go vote. Not yet! But YOU CAN! Go Vote!!! #
NYCBlackStar|instagram|0.7772|0.0|0.698|0.302|And this gif pretty much sums up the circus of an election we had! Argh! Well worth the wait to https://t.co/cHX6o7jQlY
HipstahLouis|carwash54|0.7085|0.0|0.734|0.266|"RT @carwash54: Me @ the beginning of the election: Ain't no way America letting a cheeto become president. lol what a joke Me November 7,"
himynameisjody|ImmortalTech|0.0|0.0|1.0|0.0|RT @ImmortalTech: Election night in America... https://t.co/OWC0MbDXVj
himynameisjody|twitter|0.0|0.0|1.0|0.0|RT @ImmortalTech: Election night in America... https://t.co/OWC0MbDXVj
albaugh75|ABC|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
albaugh75|abcnews|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
StanShaffer4|twitter|0.128|0.0|0.919|0.081|Was it legal for the Blk Panthers to b out for one of obamoes election in chi town? https://t.co/11uoL5g07z
mbaangluuc|DonaldJTrumpJr|-0.3595|0.098|0.902|0.0|RT @DonaldJTrumpJr: Media elites have done everything they can to stop Trump. WE THE PEOPLE will rise up and take back America! #Trump #Ele
NightlyQuest|WDFx2EU8|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
NightlyQuest|t|-0.7284|0.242|0.758|0.0|RT @WDFx2EU8: ELECTION FRAUD: Utah Election In Shambles! Democrats In Vote-By-Mail State Received Multiple Mail-In Ballots! https://t.co/7h
mouton_n0ir|twitter|0.4926|0.0|0.715|0.285|:'3some good election nite listening! get on it https://t.co/PPPkaJcYNi
jnee_roberts|mike_pence|0.0|0.0|1.0|0.0|"RT @mike_pence: This Election Day, America is standing at the crossroads of history. RT this if you're voting for @realDonaldTrump. Togethe"
mirdiy95|twitter|0.5106|0.0|0.752|0.248|If we are all being honest about tonight's election coverage...  https://t.co/KBI5mJXdWc
SDTokadam|youtube|0.0|0.0|1.0|0.0|The Young Turks Election Day Coverage 2016 https://t.co/pbqfth227U halk tvden sect take edercesine the young turks
tamaravh|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
tamaravh|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
JB93621|ABC|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
JB93621|abcnews|0.0|0.0|1.0|0.0|RT @ABC: Cake bust of Donald Trump wheeled into Trump Tower. The cake's baker said it took 50 hours to make. https://t.co/uLT42fdPGw #Elect
bustosrudy92|twitter|-0.2716|0.202|0.656|0.142|Clear example of what this election has done to this country. Utterly disgusted. https://t.co/5dXcUcwEjQ
Kat_Block_|Things4WhitePpl|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
Kat_Block_|twitter|0.0|0.0|1.0|0.0|RT @Things4WhitePpl: Breaking up over an election. https://t.co/2K3zfhewRY
MaggieBourbon|Michael_Flores|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
MaggieBourbon|rainmandigitalmedia|0.4019|0.0|0.816|0.184|RT @Michael_Flores: The #RainManShow Tainted Election special is live. #electionday #taintedelection https://t.co/SsREbMZQ7Z https://t.co/
TuNaLdO|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
TuNaLdO|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
Allison15Brandi|dansvllivan|0.9136|0.0|0.568|0.432|"RT @dansvllivan: all jokes aside, i just hope that whoever wins this election restores our country and makes it better than it already is."
Kittie0ber1968|YouTube|0.4404|0.0|0.769|0.231|I liked a @YouTube video https://t.co/hn8pMYZn6E Live Election Updates &amp; Issues That Matter | The Peoples Playhouse | 2016
Kittie0ber1968|youtube|0.4404|0.0|0.769|0.231|I liked a @YouTube video https://t.co/hn8pMYZn6E Live Election Updates &amp; Issues That Matter | The Peoples Playhouse | 2016
Shuk_bi|twitter|-0.5574|0.213|0.787|0.0|Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/7iCnZDMwBh
salemramsnj||0.0|0.0|1.0|0.0|"I posted 11 photos on Facebook in the album ""Election Day 2016 @ Salem High School"" https://t.co/tHlXt1bCfy"
salemramsnj|facebook|0.0|0.0|1.0|0.0|"I posted 11 photos on Facebook in the album ""Election Day 2016 @ Salem High School"" https://t.co/tHlXt1bCfy"
Coach_Schmitt1|twitter|0.3612|0.0|0.706|0.294|Election returns had me like #ElectionNight https://t.co/YfJTVlRncO
MamaBearTo2|twitter|0.0|0.0|1.0|0.0|Michigan Republican law makers VOTE FOR TRUMP or next election I will NOT be voting for you. 16 Electoral votes Nee https://t.co/sPn4sTdUxn
CarolCcsee|MaryLoveUS4|0.4939|0.0|0.833|0.167|RT @MaryLoveUS4: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/br0QOB4q2R https://t
CarolCcsee|thegatewaypundit|0.4939|0.0|0.833|0.167|RT @MaryLoveUS4: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/br0QOB4q2R https://t
iKendrick61|Capitals|0.0|0.0|1.0|0.0|RT @Capitals: 1 RT = 1 Vote! #VoteWilson #CapsElectionNightFollow along all day here: https://t.co/LEHLr7m9fB https://t.co/03x2pavnIz
iKendrick61|nhl|0.0|0.0|1.0|0.0|RT @Capitals: 1 RT = 1 Vote! #VoteWilson #CapsElectionNightFollow along all day here: https://t.co/LEHLr7m9fB https://t.co/03x2pavnIz
spencer_pdx|slmandel|0.3612|0.0|0.865|0.135|RT @slmandel: I went to CNN's election results page and so far it's looking a lot like LSU-Alabama. https://t.co/7ZFDXatxOf
spencer_pdx|twitter|0.3612|0.0|0.865|0.135|RT @slmandel: I went to CNN's election results page and so far it's looking a lot like LSU-Alabama. https://t.co/7ZFDXatxOf
crabtrem|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: This election my dad did not spend time raising $ from the billionaire elite. Instead he spent time talking to the Amer
chujo9|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
chujo9|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
diannemacevedo|lisforlex|0.3818|0.129|0.588|0.282|"RT @lisforlex: No matter who wins the election, Jesus will still be King "
JayceeHobbs|TexasObserver|-0.5423|0.149|0.851|0.0|RT @TexasObserver: Have you seen these dudes? @cd_hooks talks to a Fort Bend candidate who says these guys are harassing voters https://t.c
JayceeHobbs||-0.5423|0.149|0.851|0.0|RT @TexasObserver: Have you seen these dudes? @cd_hooks talks to a Fort Bend candidate who says these guys are harassing voters https://t.c
DylanWithoutBob|samsanders|0.0|0.0|1.0|0.0|RT @samsanders: Here's @NPR's live election  night blog: https://t.co/UaPBLn1Kmu
DylanWithoutBob|npr|0.0|0.0|1.0|0.0|RT @samsanders: Here's @NPR's live election  night blog: https://t.co/UaPBLn1Kmu
TXNativePatriot|bigangrylaw|0.0|0.0|1.0|0.0|"@bigangrylaw @RamonRoblesJr BTW, I am drinking beer, listening to #JimmyBuffet and grilling in the dark. What elect https://t.co/145KCLq2Me"
TXNativePatriot|twitter|0.0|0.0|1.0|0.0|"@bigangrylaw @RamonRoblesJr BTW, I am drinking beer, listening to #JimmyBuffet and grilling in the dark. What elect https://t.co/145KCLq2Me"
BlackDynamite85|CamFAwesome|0.3304|0.16|0.634|0.205|"RT @CamFAwesome: So many election parties tonight. It's going to be crazy! I hope it's ""buy a stranger a shot"" crazy, and not ""get shot by"
JenOleniczak|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
CollectedN|usatoday|0.0|0.0|1.0|0.0|News outlets preach caution on election calls https://t.co/CnHfJ2Z3JV
azcbradshaw|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
GuarimbaSiHay|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
GuarimbaSiHay|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
JasonAlt_dj|courierpostonline|0.0|0.0|1.0|0.0|"ELECTION 2016: Your one-stop place for results from Camden, Burlington &amp; Gloucester counties https://t.co/Zx5z0zEba0"
Rawadhi04|nourjafar|0.0|0.0|1.0|0.0|RT @nourjafar: I'm so afraid of the election results. https://t.co/b9yKuetFko
Rawadhi04|twitter|0.0|0.0|1.0|0.0|RT @nourjafar: I'm so afraid of the election results. https://t.co/b9yKuetFko
nelllyxo|gabbbiiieeee_|-0.8115|0.315|0.606|0.08|"RT @gabbbiiieeee_: im ready for this fucking election to be over so these racist, homophobic, ignorant ass patients in my office can shut t"
haileelovesfood|fro_zhen|-0.0772|0.226|0.557|0.217|"RT @fro_zhen: election drinking game: every state trump wins, take a shot. if he wins the election, drink until you die of alcohol poisoning"
antistuff|directv|0.0|0.0|1.0|0.0|"Check out ""Election HQ Mix"" on DIRECTV channel 347. https://t.co/4B6HeQJtcW"
deadgansey|taylorswift13|-0.1531|0.151|0.849|0.0|no shade but where has @taylorswift13 been for this election
pizdapalace|JamesOKeefeIII|0.7012|0.178|0.506|0.316|@JamesOKeefeIII is only hurting the DNC trying to RIG the election. GREAT JOB JAMES....KEEP THE TRUTH GOING!!! https://t.co/BQ10ep7z9G
pizdapalace|twitter|0.7012|0.178|0.506|0.316|@JamesOKeefeIII is only hurting the DNC trying to RIG the election. GREAT JOB JAMES....KEEP THE TRUTH GOING!!! https://t.co/BQ10ep7z9G
14Conservatives|politico|0.0|0.0|1.0|0.0|"2016 Election Results: President Live Map by State, Real-Time Voting Updates - POLITICO https://t.co/eq0vOhhSB5"
Adrienne_Young|bencasselman|0.0|0.0|1.0|0.0|RT @bencasselman: Nice.https://t.co/BUdQNjrzRE https://t.co/PLEoDcPknh
Adrienne_Young|twitter|0.0|0.0|1.0|0.0|RT @bencasselman: Nice.https://t.co/BUdQNjrzRE https://t.co/PLEoDcPknh
eruhans|biggabossben|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
eruhans|twitter|-0.3919|0.122|0.878|0.0|RT @biggabossben: When Election Day is today but you're a minority so your life was already at risk since birth https://t.co/ahbhlqkk4h
mattycakes0231|dcexaminer|0.0|0.0|1.0|0.0|RT @dcexaminer: The first polls in Florida are about to close. Full state closings and our live electoral map: https://t.co/Iz2vhOwGcW #Ele
mattycakes0231|washingtonexaminer|0.0|0.0|1.0|0.0|RT @dcexaminer: The first polls in Florida are about to close. Full state closings and our live electoral map: https://t.co/Iz2vhOwGcW #Ele
YYolanda73|electionfraud16|-0.4019|0.144|0.856|0.0|"RT @electionfraud16: Utah: Voting Machine Problems Could Force 52,000 to Use Paper Ballots - Breitbart https://t.co/iV9H8sLp7r via @Breitba"
YYolanda73|breitbart|-0.4019|0.144|0.856|0.0|"RT @electionfraud16: Utah: Voting Machine Problems Could Force 52,000 to Use Paper Ballots - Breitbart https://t.co/iV9H8sLp7r via @Breitba"
elyjiahstreeter|SavanaLuttrell|-0.7777|0.382|0.618|0.0|"RT @SavanaLuttrell: this election has me sick to my stomach, america is screwed!"
KimTroester|AlliTroester|-0.6597|0.268|0.732|0.0|"@AlliTroester gives new meaning to the election mindset of ""we're fucked either way"". "
lovedbydennis|healthandcents|-0.41|0.215|0.671|0.113|"RT @healthandcents: @payao1a1 ABSOLUTE TRUTH. If #Trump does not win this, we will never have free election again. #Globalists will control"
flatwalk|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
wcsek|PatrickMurphyFL|-0.3595|0.122|0.812|0.066|RT @PatrickMurphyFL: This is election is way too important to stay home. Lets defeat Marco Rubio -- Floridians have until 7PM to vote! #GO
SusanLenz2|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
sloepoketex|Trump2016Pence|-0.8979|0.459|0.541|0.0|"RT @Trump2016Pence: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
sloepoketex||-0.8979|0.459|0.541|0.0|"RT @Trump2016Pence: BREAKING: Florida Election Employees Caught Faking 1,000's of Stolen Absentee Ballots in Massive Voter Fraud https://t."
MirentxuCastro|washingtonpost|-0.5859|0.257|0.743|0.0|"The Fix: Donald Trump's Election Day insinuations of voter fraud, explained https://t.co/V8ZPzSxjtS"
victory1261|ChicagoDailyNew|-0.3182|0.161|0.839|0.0|RT @ChicagoDailyNew: How Write-In Ballots Could Delay Results on Election Day https://t.co/0sAXMZ4L9m https://t.co/ZXU7jBUysV
victory1261|nbcchicago|-0.3182|0.161|0.839|0.0|RT @ChicagoDailyNew: How Write-In Ballots Could Delay Results on Election Day https://t.co/0sAXMZ4L9m https://t.co/ZXU7jBUysV
Kashii_Nap|blvckpapii|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
Kashii_Nap|twitter|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
MaryJaneDaum|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
theashleymatt|LeoDiCaprio|0.0|0.0|1.0|0.0|"I know it's all about the US election tonight, but here's this again anyway. @LeoDiCaprio @NatGeo #BeforeTheFlood https://t.co/jZYgEPUAB6"
theashleymatt|channel|0.0|0.0|1.0|0.0|"I know it's all about the US election tonight, but here's this again anyway. @LeoDiCaprio @NatGeo #BeforeTheFlood https://t.co/jZYgEPUAB6"
debbiedo58|AP_Politics|0.3818|0.0|0.867|0.133|"RT @AP_Politics: On Election Day, Trump refuses to say whether he'll accept the election results. #Election2016 https://t.co/UeZzVNFgJj htt"
debbiedo58|apnews|0.3818|0.0|0.867|0.133|"RT @AP_Politics: On Election Day, Trump refuses to say whether he'll accept the election results. #Election2016 https://t.co/UeZzVNFgJj htt"
gypsybae|GAVlNREACTS|0.6249|0.0|0.661|0.339|RT @GAVlNREACTS: A great way to start Election Day https://t.co/yr6QAP3orF
gypsybae|twitter|0.6249|0.0|0.661|0.339|RT @GAVlNREACTS: A great way to start Election Day https://t.co/yr6QAP3orF
srslymikaylarae|ginapalmieri3|0.0|0.0|1.0|0.0|RT @ginapalmieri3: $1 burritos at miguel's cuz election day 
ClarissaSchreed|TheDailyShow|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
ClarissaSchreed|cc|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
JamesWilliams9|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
JamesWilliams9||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
Quinnb00b|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
Quinnb00b|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
usfreedom12|usfreedom12|0.7906|0.0|0.692|0.308|"RT @usfreedom12: @girlposts @DrMartyFox Stronger together is only good till election, after that she give u the middle finger like the Bern"
Esteban281997|nickatnyteYT|0.2023|0.0|0.913|0.087|"RT @nickatnyteYT: Got it back. Top 100 Global for the day, pushing complete.. time to tune into election night. https://t.co/ebUKnOnxCx"
Esteban281997|twitter|0.2023|0.0|0.913|0.087|"RT @nickatnyteYT: Got it back. Top 100 Global for the day, pushing complete.. time to tune into election night. https://t.co/ebUKnOnxCx"
majiktinkerbell|hockeydeb21|-0.4466|0.257|0.616|0.128|RT @hockeydeb21: LEAKED CLINTON INTERNAL DOCUMENT: Discourage Trump Supporters with Bogus Polls and Declaring Election Over https://t.co/cJ
majiktinkerbell|t|-0.4466|0.257|0.616|0.128|RT @hockeydeb21: LEAKED CLINTON INTERNAL DOCUMENT: Discourage Trump Supporters with Bogus Polls and Declaring Election Over https://t.co/cJ
CultureInStereo|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
CultureInStereo|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
Brooke_Baldwinx|kornfan_420|-0.6808|0.187|0.813|0.0|RT @kornfan_420: Was just told it's ELECTION day not ERECTION day what the hell am I supposed to do with this thing
Fleyfall|CherOfficiaI|0.6633|0.0|0.783|0.217|RT @CherOfficiaI: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
LaudyLoo|NerdylilGuy|0.0|0.0|1.0|0.0|"@NerdylilGuy listen, you made a public comment on social media about a hot topic subject, immigration...on election night. Is it really that"
Paulhardingjr|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
Heathah_|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
JehseaLynn|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
JehseaLynn|thehill|-0.5574|0.205|0.795|0.0|"RT @thehill: 2 election clerks fired in Florida for not following ""procedure and policy"" https://t.co/UQs4nrMwsr https://t.co/RIY1YMSaCc"
Eren_360|hannah_whit23|0.5719|0.0|0.709|0.291|RT @hannah_whit23: Happy Election Day to all you dreamers https://t.co/ldpJtNKFg1
Eren_360|twitter|0.5719|0.0|0.709|0.291|RT @hannah_whit23: Happy Election Day to all you dreamers https://t.co/ldpJtNKFg1
SheilaChilds1|StatesPoll|0.0|0.0|1.0|0.0|"RT @StatesPoll: My Prediction of #Election2016 11/07/2016(Final)More Details, Read my post: https://t.co/oExiU0xTRc#TrumpTrain #Trump2016"
SheilaChilds1|statespoll|0.0|0.0|1.0|0.0|"RT @StatesPoll: My Prediction of #Election2016 11/07/2016(Final)More Details, Read my post: https://t.co/oExiU0xTRc#TrumpTrain #Trump2016"
everafterwelive|anhz00|0.4574|0.0|0.857|0.143|@anhz00 @snee_jpg @maddiecarina many democrats are voting third party this election is what i (and i think maddie too) am saying!
karlyn_darlin|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
karlyn_darlin|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
breebacon20|google|0.0|0.0|1.0|0.0|My browser is going to stay on the @google election results page all night.
1Thunder_Struck|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
1Thunder_Struck|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
____Cilla|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
____Cilla|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
CamaroKiddos|DonaldJTrumpJr|0.5574|0.0|0.777|0.223|RT @DonaldJTrumpJr: Early indications: twice as many voters want a strong leader this election than in 2012. #MAGA #ElectionDay
efairhurst|fortune|-0.4588|0.25|0.75|0.0|Mean Girls Fans Are Arguing About Their Own Election https://t.co/ey8cX4taXF
WeirMB|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
WeirMB|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
mirrormatt86|channeltennews|-0.7906|0.318|0.682|0.0|"RT @channeltennews: UPDATE: @LAtimes report 1 person is dead, multiple injured following shooting near polling station. #Electionday   http"
StephCornellier|theScore|0.0|0.0|1.0|0.0|RT @theScore: VIDEO: The @Capitals are holding a bobblehead vote on U.S. #ElectionNight. https://t.co/ObRLda8xmX https://t.co/ZSkGldSFDn
StephCornellier|thescore|0.0|0.0|1.0|0.0|RT @theScore: VIDEO: The @Capitals are holding a bobblehead vote on U.S. #ElectionNight. https://t.co/ObRLda8xmX https://t.co/ZSkGldSFDn
BernardRadcliff|Rosenchild|0.0258|0.0|0.945|0.055|"RT @Rosenchild: U.S., British and German Officials say Russia's interference in the Election and backing of Trump are Unprecedented https:/"
BernardRadcliff||0.0258|0.0|0.945|0.055|"RT @Rosenchild: U.S., British and German Officials say Russia's interference in the Election and backing of Trump are Unprecedented https:/"
SgtMelons|HRC4Prison|-0.6908|0.228|0.722|0.049|"RT @HRC4Prison: DISTRACTIONWhile media tries to focus your attention on this, they want to distract you from election fraud &amp; Clinton th"
mommom_dayton|washingtonpost|0.0|0.0|1.0|0.0|Russian TV is showing nude Melania Trump and election rigging ahead of U.S. election https://t.co/xm4bAvRQ51
nomandatesDKos|nomandatesDKos|0.0|0.0|1.0|0.0|RT @nomandatesDKos: .@RepZoeLofgren: @RepMikeHonda deserves re-election to Congress in #ca17 https://t.co/EZ7FycdljC @mikehonda17
nomandatesDKos|mercurynews|0.0|0.0|1.0|0.0|RT @nomandatesDKos: .@RepZoeLofgren: @RepMikeHonda deserves re-election to Congress in #ca17 https://t.co/EZ7FycdljC @mikehonda17
katerbrts|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
katerbrts|google|0.0|0.0|1.0|0.0|RT @google: See #ElectionDay results unfold in real time on Google Search  https://t.co/dKfOxCFm2m https://t.co/CnCrDxVEfq
dejean76|Rach_IC|0.4939|0.0|0.833|0.167|RT @Rach_IC: Ugh... More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/R0yTMEIzBb
dejean76|thegatewaypundit|0.4939|0.0|0.833|0.167|RT @Rach_IC: Ugh... More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/R0yTMEIzBb
LyndaKelly|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
LyndaKelly|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
AshamedNot|Vendetta92429|0.6588|0.0|0.672|0.328|RT @Vendetta92429: Off to a great start in New Hampshire!#ElectionNight#TrumpTriumphhttps://t.co/z7GP1ueggp https://t.co/khQR80m183
AshamedNot|twitter|0.6588|0.0|0.672|0.328|RT @Vendetta92429: Off to a great start in New Hampshire!#ElectionNight#TrumpTriumphhttps://t.co/z7GP1ueggp https://t.co/khQR80m183
ShanaTargosz|twitter|0.6369|0.0|0.704|0.296|This is the best election day tweet I've seen today. https://t.co/5XT54DcEOf
BenMoull|toddpruzan|-0.3802|0.11|0.89|0.0|RT @toddpruzan: Seemed odd Trump books his election-night wake at the Hilton. Why give away the business? Until I realized! He's going to s
CruisingWes|DrJosephWarren|0.6369|0.0|0.741|0.259|Take a walk through history on the Freedom Trail for Election Day.https://t.co/IYummseRcl @DrJosephWarren https://t.co/Rl8f7WQeTy
CruisingWes|twitter|0.6369|0.0|0.741|0.259|Take a walk through history on the Freedom Trail for Election Day.https://t.co/IYummseRcl @DrJosephWarren https://t.co/Rl8f7WQeTy
MichaelDupuis4|DonaldJTrumpJr|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you VOTED TO DRAIN THE SWAMP! #MAGA #ElectionDay #Election https://t.co/TkUPGBNYkg
MichaelDupuis4|twitter|0.0|0.0|1.0|0.0|RT @DonaldJTrumpJr: RT if you VOTED TO DRAIN THE SWAMP! #MAGA #ElectionDay #Election https://t.co/TkUPGBNYkg
valley0fwolves|Terravitabass|0.5093|0.0|0.829|0.171|RT @Terravitabass: Got to vote on weed and porn in the election today. Welcome to California! https://t.co/9UnmX9AaJ1
valley0fwolves|twitter|0.5093|0.0|0.829|0.171|RT @Terravitabass: Got to vote on weed and porn in the election today. Welcome to California! https://t.co/9UnmX9AaJ1
1stThunderThief|hrtablaze|0.9207|0.0|0.645|0.355|RT @hrtablaze: My Bernie Sanders loving nephew who has been messing with me all election just told me he voted TRUMP !!! WOOT WOOT ! #elect
siaayrom|FrankLuntz|0.4019|0.0|0.891|0.109|"RT @FrankLuntz: All eyes will be in Virginia for 2017.Tim Kaine's Senate seat will open up, and they will have a special election.  #Elec"
DerrickMinor|twitter|-0.2263|0.112|0.888|0.0|These two are anxiously awaiting the election results. Especially the one on the right. #Election2016 https://t.co/jBpdmoeZMI
frazier_ann|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
GCC_legal|reuters|-0.4404|0.209|0.791|0.0|RT ReutersOpinion: The psychology behind voters' choices  and election madness: https://t.co/8zq9jn04Xu https://t.co/EXYhCfBsQ3
MSMuralles|SenSanders|0.6705|0.0|0.744|0.256|RT @SenSanders: Election Day should be a national holiday so that everyone has the time and opportunity to vote.
jeshizaemon|fivethirtyeight|-0.0173|0.215|0.574|0.211|This is awful. Poling Place shooting in Azusa D: https://t.co/80vhjyaCAq
ortizylime|Evil_Dumbledore|-0.6486|0.212|0.677|0.111|"RT @Evil_Dumbledore: Can't wait until this election is over so we can go back to hating each other for shit that matters, like ford vs chev"
mikethemoody|digitalrailgun|0.4199|0.0|0.843|0.157|RT @digitalrailgun: Ready for the election here in Vancouver! @TYTPolitics @TYTNetwork @cenkuygur @JordanChariton #TYT #tytlive #ElectionDa
donkler|YouTube|0.4753|0.0|0.808|0.192|I liked a @YouTube video from @scrowder https://t.co/QZbdNSNi1O Crowder's ALL-STAR Election Live Stream! | Louder With Crowder
donkler|youtube|0.4753|0.0|0.808|0.192|I liked a @YouTube video from @scrowder https://t.co/QZbdNSNi1O Crowder's ALL-STAR Election Live Stream! | Louder With Crowder
yurbaink|cnni|0.6369|0.0|0.833|0.167|"RT @cnni: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/0RU6ozSJGg"
yurbaink|cnn|0.6369|0.0|0.833|0.167|"RT @cnni: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/0RU6ozSJGg"
jNaemaraj|MASEEZUSWEST|0.0|0.0|1.0|0.0|RT @MASEEZUSWEST: The election effects the whole world soo https://t.co/EcG4osFmCI
jNaemaraj|twitter|0.0|0.0|1.0|0.0|RT @MASEEZUSWEST: The election effects the whole world soo https://t.co/EcG4osFmCI
LeAnne_Stokes|OANN|0.0|0.0|1.0|0.0|RT @OANN: All hands on deck at #OANN today! Election Day coverage starts in just under 30 minutes (7 PM EST)! #TuneIn for the latest from t
TrumpWithUSA|carrieksada|0.7964|0.0|0.664|0.336|RT @carrieksada: Please listen to the remarkable @LouDobbs as he shares what is at stake in this election:#MAGA https://t.co/I5djUZ8CVJ
TrumpWithUSA|twitter|0.7964|0.0|0.664|0.336|RT @carrieksada: Please listen to the remarkable @LouDobbs as he shares what is at stake in this election:#MAGA https://t.co/I5djUZ8CVJ
Heidic282|rascalblog|0.0258|0.158|0.712|0.13|RT @rascalblog: I bloody love US election nights. But this is the first one where I've been worried about what the result will do to the Do
MadridMagical|MJosephSheppard|0.7506|0.0|0.701|0.299|RT @MJosephSheppard: Pinellas County Florida Obama won by 5.6 Current two party vote GOP 55% Dem 45%https://t.co/G1z7oNy6Yf
MadridMagical|votepinellas|0.7506|0.0|0.701|0.299|RT @MJosephSheppard: Pinellas County Florida Obama won by 5.6 Current two party vote GOP 55% Dem 45%https://t.co/G1z7oNy6Yf
EltonAJMenezes|ABCWorldNews|0.4019|0.0|0.881|0.119|RT @ABCWorldNews: TUNE-IN: Special election night edition of #WorldNewsTonight is live on the east coast right now - RT if you're watching
TheRealWize|lsarsour|0.8479|0.0|0.638|0.362|"RT @lsarsour: I hope that if this election taught Muslim Americans anything, is that's it more important to be respected than accepted. #My"
Eddie_Here|IMPaulWilliams|0.6428|0.065|0.695|0.239|RT @IMPaulWilliams: Heading for London and the @ASCAP London Awards. Missing the election news but I voted.  Life is good.   https://t.
Eddie_Here||0.6428|0.065|0.695|0.239|RT @IMPaulWilliams: Heading for London and the @ASCAP London Awards. Missing the election news but I voted.  Life is good.   https://t.
Laia_QR|nytimes|0.0|0.0|1.0|0.0|Presidential Election Results https://t.co/4gIu05Kec1
mikemcfillin|InappropriateSB|0.0|0.0|1.0|0.0|RT @InappropriateSB: This election in a nutshell https://t.co/TE1m8Scmmi
mikemcfillin|twitter|0.0|0.0|1.0|0.0|RT @InappropriateSB: This election in a nutshell https://t.co/TE1m8Scmmi
Adhirizkyputra|AJEnglish|0.0|0.0|1.0|0.0|RT @AJEnglish: Here's when to expect election results.Follow the live results here: https://t.co/arXvIMQVja #ElectiondDay #Election2016 ht
Adhirizkyputra|interactive|0.0|0.0|1.0|0.0|RT @AJEnglish: Here's when to expect election results.Follow the live results here: https://t.co/arXvIMQVja #ElectiondDay #Election2016 ht
sophieissoapy|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
sophieissoapy|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
JohnnyT2413|MikeDrucker|0.4404|0.0|0.888|0.112|"RT @MikeDrucker: If you have time today, go back and watch some of @LateNightSeth's closer look segments and witness how good he's been thi"
NCNShelenberger|twitter|0.0|0.0|1.0|0.0|A 33-year-old man explains why  this election prompted him to vote for the first time. #PAelectionCNHI https://t.co/sZXW0Ajs4x
finallyzach|aqxurs|0.0|0.0|1.0|0.0|@aqxurs also there has never been a case in history where a rogue electoral college member has changed the result of an election
aliciachavez_3|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
syaldram|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
kiki_designs|annehelen|0.6369|0.0|0.811|0.189|.@annehelen @maramcewin I love how telling the one way signs are... in this election...only one way to go #ImWithHer  @HillaryClinton
BeingFarhad|twitter|-0.5574|0.195|0.805|0.0|RT Donald Trump keeps telling us that the election is rigged. So what's the real risk of #voterfraud today? https://t.co/JbI3VkTAo7 #f4f #
sumonszzd|mashable|0.0|0.0|1.0|0.0|America gets lit: The Lite Brite guide to election results https://t.co/TSWscJJ9Tb
lucie_harris|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
lucie_harris|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: How other countries would vote in the American election https://t.co/kYiIOsGYO0 https://t.co/eoQw7s3H8V
corellianjedi2|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
corellianjedi2|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
evanway|SidneyCrosbyEgo|0.765|0.0|0.752|0.248|RT @SidneyCrosbyEgo: The best part about election day is that we get to watch McDavid and Crosby play before the world ends.
ayeejanae|kayyebby|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
ayeejanae|twitter|0.5994|0.0|0.794|0.206|RT @kayyebby: your wcw thinks election day &amp; inauguration day are the same thing lmao https://t.co/V1aloSIhj0
ThomasAHester2|spkhp|0.4588|0.0|0.833|0.167|RT @spkhp: Here's a thread of quotes from my kids about Election Day. In case anyone cares.
kf4bef|WalidPhares|0.0|0.0|1.0|0.0|RT @WalidPhares: Follow returns and results here https://t.co/I6vf12RUIk
kf4bef|foxnews|0.0|0.0|1.0|0.0|RT @WalidPhares: Follow returns and results here https://t.co/I6vf12RUIk
lizthemermaid|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
lizthemermaid||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
BeckermanJosh|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
BeckermanJosh|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
stephenjstedman|eosnos|0.3612|0.0|0.898|0.102|"RT @eosnos: ""Looking at exit polls is like hooking up with your ex-girlfriend. You know before you do it that you shouldnt."" https://t.co/"
stephenjstedman|t|0.3612|0.0|0.898|0.102|"RT @eosnos: ""Looking at exit polls is like hooking up with your ex-girlfriend. You know before you do it that you shouldnt."" https://t.co/"
_jcm11|immigrant4trump|0.7506|0.0|0.766|0.234|"RT @immigrant4trump: If you make this go viral, Trump will win. It's about 2 minutes that makes the choice in this election crystal clear h"
Zipfireteam|mashable|0.0|0.0|1.0|0.0|Australia offers 'democracy sausages' to Americans in their hour of need- Don't wo https://t.co/ch2qUfJOwH
FewerHorsesNBay|MakeupArtistmag|0.0|0.0|1.0|0.0|RT @MakeupArtistmag: We're voting for the 'SNL' make-up/hair team for their Hillary Clinton and Donald Trump transformations! https://t.co/
FewerHorsesNBay|t|0.0|0.0|1.0|0.0|RT @MakeupArtistmag: We're voting for the 'SNL' make-up/hair team for their Hillary Clinton and Donald Trump transformations! https://t.co/
9ineWaves|heybri_|0.0|0.0|1.0|0.0|RT @heybri_: *pours coconut oil on this election*
BreezyBiz|JeffProbst|0.0|0.0|1.0|0.0|Hey @JeffProbst how long do you think it'll take you to read all of the election votes Survivor-style?
ladiharli|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
listelian|land_planarian|0.2023|0.0|0.859|0.141|RT @land_planarian: Erowid Sarah Palin's election coverage has been top notch https://t.co/TiHwjMQGHA
listelian|twitter|0.2023|0.0|0.859|0.141|RT @land_planarian: Erowid Sarah Palin's election coverage has been top notch https://t.co/TiHwjMQGHA
LeahLikesDogs|vcrichardson|0.0|0.0|1.0|0.0|@vcrichardson when the stakes aren't as high as for election cupcakes
StephCavazos14|AC360|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
StephCavazos14|t|0.743|0.105|0.576|0.319|"RT @AC360: .@ananavarro: ""It would be sweet, sweet justice if tonight it was the Latino vote that defeated Donald Trump"" https://t.co/ZTdYJ"
dagraffman|dsudis|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
dagraffman|twitter|0.7772|0.0|0.639|0.361|RT @dsudis: Ida B. Wells getting the love on Election Day in Chicago!! https://t.co/GGG2p4sV43
CDaudette|THE_KURZE|-0.7909|0.25|0.75|0.0|@THE_KURZE so many people don't understand their votes mean nothing. I hope this election has shown people that our gov is corrupt as hell.
PharaohJ7|TheOnion|0.0|0.0|1.0|0.0|"RT @TheOnion: Presenting our Election Day live blog, bringing readers up-to-the-minute coverage they neither asked for nor deserve https://"
PharaohJ7||0.0|0.0|1.0|0.0|"RT @TheOnion: Presenting our Election Day live blog, bringing readers up-to-the-minute coverage they neither asked for nor deserve https://"
SunnyJL52|EricTrump|0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
SunnyJL52||0.5562|0.0|0.86|0.14|"RT @EricTrump: On the eve of this election, let's always remember our bravest men &amp; women who sacrificed everything for our nation! https:/"
misstozak|jerome_corsi|-0.5859|0.153|0.847|0.0|RT @jerome_corsi: TRUMP NEEDS ALL POSSIBLE VOTERS IN PA - voter fraud being reported EVENING HOURS WILL DECIDE ELECTION - get all Trump vot
boodygoon|JelvinParra13|0.0|0.0|1.0|0.0|RT @JelvinParra13: These are the recent polls of the presidential election: https://t.co/MtZWdfYwKT
boodygoon|twitter|0.0|0.0|1.0|0.0|RT @JelvinParra13: These are the recent polls of the presidential election: https://t.co/MtZWdfYwKT
LoliLoli2823|AllenWest|0.0|0.0|1.0|0.0|RT @AllenWest: I'll be on CBS DFW live. Election coverage starts at 6pm CT with updates twice each hour. Watch it streaming here: https://t
LoliLoli2823||0.0|0.0|1.0|0.0|RT @AllenWest: I'll be on CBS DFW live. Election coverage starts at 6pm CT with updates twice each hour. Watch it streaming here: https://t
AccessSanDiego|10news|0.6467|0.0|0.808|0.192|"Happy election day ""I VOTED!"" sticker gives you these deals! Election Day Deals: Doughnuts and Uber rides -... https://t.co/XMLjlITILO"
a_perrrr|lpdanoodlehead|-0.6124|0.4|0.6|0.0|RT @lpdanoodlehead: I'm terrified about this election.
GCC_legal|reuters|0.0|0.0|1.0|0.0|RT ReutersPolitics: Factbox: State-by-state poll closing times for U.S. election https://t.co/ykuKzUBo4Z https://t.co/0aV13wVq9Z
caramelambition|illpatic|0.5719|0.0|0.802|0.198|RT @illpatic: The new North Carolina state flag if Gov. McCrory wins re-election tonight #FlyTheL https://t.co/Kq4r42HCAJ
caramelambition|twitter|0.5719|0.0|0.802|0.198|RT @illpatic: The new North Carolina state flag if Gov. McCrory wins re-election tonight #FlyTheL https://t.co/Kq4r42HCAJ
Darksbane7|CNN|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
Darksbane7|twitter|-0.2732|0.084|0.875|0.042|"RT @CNN: Its all up to you now. No matter who youre voting for, see your vote counted on CNN election night in America.  https://t.co/8"
christylynn923|isardasorensen|0.0|0.0|1.0|0.0|"RT @isardasorensen: The @EmpireStateBldg shines red, white &amp; blue on this historic #ElectionNight in America. #election #ElectionDay  #NYC"
GateKeeper1776|healthandcents|-0.41|0.215|0.671|0.113|"RT @healthandcents: @payao1a1 ABSOLUTE TRUTH. If #Trump does not win this, we will never have free election again. #Globalists will control"
ManitobaRetweet|BrittAtGlobal|0.0|0.0|1.0|0.0|RT @BrittAtGlobal: Plan on viewing #USElection2016 tonight? Here's a list of places around #Winnipeg to watch https://t.co/px4ozgJqX8
ManitobaRetweet|globalnews|0.0|0.0|1.0|0.0|RT @BrittAtGlobal: Plan on viewing #USElection2016 tonight? Here's a list of places around #Winnipeg to watch https://t.co/px4ozgJqX8
GeorgiaDaskalos|DRUDGE_REPORT|0.3182|0.0|0.827|0.173|RT @DRUDGE_REPORT: Madonna breaks promise to give oral to Hillary voters... https://t.co/obsQ3RlTFO
GeorgiaDaskalos|nydailynews|0.3182|0.0|0.827|0.173|RT @DRUDGE_REPORT: Madonna breaks promise to give oral to Hillary voters... https://t.co/obsQ3RlTFO
mskerryd|nicole|0.4019|0.0|0.816|0.184|@nicole I just inhaled half the chips I was bringing to my friend's Election party. 
JonaPrelvukaj|deadmau5|0.0|0.0|1.0|0.0|RT @deadmau5: Election night starter kit: https://t.co/eWLzxyPhQ3
JonaPrelvukaj|twitter|0.0|0.0|1.0|0.0|RT @deadmau5: Election night starter kit: https://t.co/eWLzxyPhQ3
skorpyos|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
skorpyos|politico|0.0|0.0|1.0|0.0|RT @politico: Polls are about to close in multiple states. Follow live results here: https://t.co/YYB0l0V0BN https://t.co/lW4cC0Gvaj
joannele2001|ForTrump|0.3182|0.0|0.909|0.091|RT @ForTrump: Please get out and vote. Do not listen 2exit polls. This is the election that will decide our country's future.  Let's #MAGA
ggindc|ABCPolitics|0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
ggindc||0.0|0.0|1.0|0.0|"RT @ABCPolitics: NEW: Nearly 7 in 10 North Carolina voters oppose HB2, the so-called ""bathroom bill,"" per preliminary exit polls https://t."
Augied5|twitter|0.3612|0.0|0.615|0.385|Watching the election like https://t.co/kATbY1kTNF
RabNelzan|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
RabNelzan|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
TheAFactor15|SoaRPraizist|0.5719|0.0|0.802|0.198|"RT @SoaRPraizist: If Trump wins the election, I will make artwork for everyone that RTs this tweet"
Colak|AnsonWhaley|0.0|0.0|1.0|0.0|RT @AnsonWhaley: This is absolutely the only way the first vote could have been registered in this election. https://t.co/qhoJ4AJe0q
Colak|vine|0.0|0.0|1.0|0.0|RT @AnsonWhaley: This is absolutely the only way the first vote could have been registered in this election. https://t.co/qhoJ4AJe0q
renukamendiss|JohnIbbitson|0.0|0.0|1.0|0.0|RT @JohnIbbitson: I just sent in my contribution to an election pool. Somehow I feel obligated to go on the record. So:Clinton: 329 ecvTr
Sundip|NateSilver538|0.0|0.0|1.0|0.0|RT @NateSilver538: So here's the link to our election night model! Forecast will update as states are CALLED (not on partial returns): http
WNYC|wnyc|0.0|0.0|1.0|0.0|"As #ElectionNight results come in, WNYC will have the latest right here: https://t.co/EJuQ41zVER https://t.co/RM4ObRf99g"
khcopeland1|JoeBiden|0.0|0.0|1.0|0.0|RT @JoeBiden: There are world-class candidates running at all levels in this election. Vote down the line for Democrats who will keep us mo
ootdyo|MTVNews|0.0|0.0|1.0|0.0|RT @MTVNews: our livestream is starting. we've got @JulianneRoss and @GabyWilson chopping it up about the election with @PUSHA_T! https://t
ootdyo||0.0|0.0|1.0|0.0|RT @MTVNews: our livestream is starting. we've got @JulianneRoss and @GabyWilson chopping it up about the election with @PUSHA_T! https://t
AREEV1|HipHopzilla|0.0|0.0|1.0|0.0|RT @HipHopzilla: Colin Kaepernick Says He Won't Vote in 2016 Presidential Election https://t.co/5YSxaJdeL9
AREEV1|hiphopzilla|0.0|0.0|1.0|0.0|RT @HipHopzilla: Colin Kaepernick Says He Won't Vote in 2016 Presidential Election https://t.co/5YSxaJdeL9
Deruelle20_|SidneyCrosbyEgo|0.765|0.0|0.752|0.248|RT @SidneyCrosbyEgo: The best part about election day is that we get to watch McDavid and Crosby play before the world ends.
jasmynph0|burgurll|0.0|0.0|1.0|0.0|"RT @burgurll: Michellle Obama should run for president next election and her slogan should be ""Ya'll thought we were done"""
PattiDudek|rjcc|0.0|0.0|1.0|0.0|"RT @rjcc: Another trend to follow is the hashtag #CripTheVote, tracking the experiences of people with disabilities voting. https://t.co/RQ"
PattiDudek|t|0.0|0.0|1.0|0.0|"RT @rjcc: Another trend to follow is the hashtag #CripTheVote, tracking the experiences of people with disabilities voting. https://t.co/RQ"
laurnorman|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
laurnorman|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
LaurenIsTheBoss|AllyBrooke|0.7506|0.0|0.575|0.425|RT @AllyBrooke: Praying for our election tomorrow and may God bless our country 
JMawhirter|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
JMawhirter|businessinsider|0.5719|0.0|0.821|0.179|RT @businessinsider: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/E3uNuK6fMw https://t.c
SantoFanara|IZOD|0.296|0.0|0.833|0.167|RT @IZOD: America votes. Join the Election Day conversation with #MyVote2016 https://t.co/BWuiwAxas6
SantoFanara|twitter|0.296|0.0|0.833|0.167|RT @IZOD: America votes. Join the Election Day conversation with #MyVote2016 https://t.co/BWuiwAxas6
bad_indian_girl|Milbank|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
bad_indian_girl|twitter|0.3612|0.06|0.815|0.124|RT @Milbank: They built a cash bar at Trump election night party-- and his supporters are going to pay for it. https://t.co/X18u0HieSN
nehapatel620|twitter|-0.4767|0.119|0.881|0.0|I know I've been spamming with election tweets  But here is my final 1 before we all find out b/c it was my 1st ti https://t.co/wNIymZ3zGq
c_thegerg|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
c_thegerg|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
SicilianIrish02|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Donald #Trump. Follow @nbcconnecticut for the latest election news.https://t.co/S7TjIfwe65
celesteka|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
Eric__TH|VoiceOverDan|0.6801|0.0|0.741|0.259|RT @VoiceOverDan: I'm really hoping this election night ends up being like game 5 against the Thunder in 2012.
mlafferty1|CaitlinDineen|0.296|0.0|0.879|0.121|@CaitlinDineen Here's yer election night pizza at the Villages Daily Sun. I'm helping edit there tonight. https://t.co/JaUXrMAQXs
mlafferty1|twitter|0.296|0.0|0.879|0.121|@CaitlinDineen Here's yer election night pizza at the Villages Daily Sun. I'm helping edit there tonight. https://t.co/JaUXrMAQXs
taytayheyhey_|kimberly_carden|0.0|0.0|1.0|0.0|"RT @kimberly_carden: people ask why i'm not as concerned about the election as i ""should"" be https://t.co/SpGgMg2yBV"
taytayheyhey_|twitter|0.0|0.0|1.0|0.0|"RT @kimberly_carden: people ask why i'm not as concerned about the election as i ""should"" be https://t.co/SpGgMg2yBV"
randypittman71|NBCNews|0.0|0.0|1.0|0.0|"RT @NBCNews: It's just minutes until polls close in Georgia, Indiana, Kentucky, South Carolina, Vermont &amp; Virginia. Follow here: https://t."
randypittman71||0.0|0.0|1.0|0.0|"RT @NBCNews: It's just minutes until polls close in Georgia, Indiana, Kentucky, South Carolina, Vermont &amp; Virginia. Follow here: https://t."
AshleyRaulet|WFTV|0.0|0.0|1.0|0.0|RT @WFTV: #Election results are beginning to come in: https://t.co/01VQr3a43C
AshleyRaulet|wftv|0.0|0.0|1.0|0.0|RT @WFTV: #Election results are beginning to come in: https://t.co/01VQr3a43C
JaniceR09496229|janeosanders|0.6369|0.071|0.66|0.269|"RT @janeosanders: Nice story &amp; video re: our incredible supporters  tough day, various choices. #OurRevolution endures. https://t.co/E6Vbi"
JaniceR09496229|t|0.6369|0.071|0.66|0.269|"RT @janeosanders: Nice story &amp; video re: our incredible supporters  tough day, various choices. #OurRevolution endures. https://t.co/E6Vbi"
ToniStinchcomb|SarahWoodwriter|0.0|0.0|1.0|0.0|RT @SarahWoodwriter: Sometimes you just need to dance with your dogs to Bob Marley to prepare yourself for Election Day.  https://t.co/
ToniStinchcomb|t|0.0|0.0|1.0|0.0|RT @SarahWoodwriter: Sometimes you just need to dance with your dogs to Bob Marley to prepare yourself for Election Day.  https://t.co/
wmsal7|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
marinaslater|parleyxxx|0.0516|0.202|0.588|0.21|RT @parleyxxx: To ease election day anxiety: #marinelife suspended in light and time in their natural environment. https://t.co/X69RwX4ZuZ
marinaslater|parley|0.0516|0.202|0.588|0.21|RT @parleyxxx: To ease election day anxiety: #marinelife suspended in light and time in their natural environment. https://t.co/X69RwX4ZuZ
candynheba|ladygaga|0.0|0.0|1.0|0.0|RT @ladygaga: RT and spread this message Monsters! It's election KRUNCHTime and EVERY VOTE counts! #ElectionDay #Elections2016 #GoVote #Vot
aalanadelreyy|diego_goes_|0.0|0.0|1.0|0.0|"RT @diego_goes_: Election Day go out and vote, unless you're voting for trump then that's tomorrow"
superfabis|theverge|0.0|0.0|1.0|0.0|10 provocative political novels to read after the election https://t.co/4jIz30so5N https://t.co/VA6nLII59q
tinyceli_|KathleenLights1|0.4199|0.141|0.573|0.286|RT @KathleenLights1: Hope everyone voted today! This election has traumatized me.... I pray for America.
whatmsees|HIGH_TIMES_Mag|0.2225|0.0|0.921|0.079|RT @HIGH_TIMES_Mag: We're back on FB Live! Want to know the second weed gets legalized? IGH TIMES is covering the election live! https://t.
whatmsees||0.2225|0.0|0.921|0.079|RT @HIGH_TIMES_Mag: We're back on FB Live! Want to know the second weed gets legalized? IGH TIMES is covering the election live! https://t.
blessed4home|realDonaldTrump|0.7836|0.0|0.723|0.277|RT @realDonaldTrump: I will be watching the election results from Trump Tower in Manhattan with my family and friends. Very exciting!
kimwhocries|TheLastRefuge2|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
kimwhocries|twitter|-0.4588|0.214|0.786|0.0|"RT @TheLastRefuge2: Typical Nevada Politics.  Election Officials/Workers wearing ""Defeat Trump"" T-Shirts. https://t.co/TqlBqmjy0G"
elmorephd|MissD4Trump|-0.4738|0.123|0.877|0.0|RT @MissD4Trump: This election will be decided by the people working 2 to 3 jobs.We need your vote! We need your evening vote! Ignore the T
SunnyAtTheGulf|IngrahamAngle|0.0|0.0|1.0|0.0|"RT @IngrahamAngle: Will Obama's ""election monitors"" do anything about this?? https://t.co/oMpf1nimAQ"
SunnyAtTheGulf|twitter|0.0|0.0|1.0|0.0|"RT @IngrahamAngle: Will Obama's ""election monitors"" do anything about this?? https://t.co/oMpf1nimAQ"
CurrentSocials|mashable|0.0|0.0|1.0|0.0|#SM America gets lit: The Lite Brite guide to election results: The 2016 presidential https://t.co/DgQM4A9tN9
hey_its_bai|PaperWash|0.3612|0.0|0.878|0.122|RT @PaperWash: Here is what the electoral map would look like if only bakers voted in the election https://t.co/Y0w3utclBq
hey_its_bai|twitter|0.3612|0.0|0.878|0.122|RT @PaperWash: Here is what the electoral map would look like if only bakers voted in the election https://t.co/Y0w3utclBq
BlueEyedRobin|youtube|0.0|0.0|1.0|0.0|Keeping up election year traditions https://t.co/kTqI5eyZSn #mydatewiththepresidentsdaughter
suidfc|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/FbSc1sQ8jN
suidfc|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/FbSc1sQ8jN
ryanpitts|mattdennewitz|0.0|0.0|1.0|0.0|@mattdennewitz what does Pitchfork eat on election night?
SluttyVanessaC|xvideos|-0.8553|0.54|0.46|0.0|Tired of this election bullshit?  Jerk off to my videos instead!https://t.co/i2E1FvbtwM
orataiculhane|LeahR77|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
orataiculhane|breitbart|0.8061|0.0|0.673|0.327|RT @LeahR77: Exits! Exits! Exits! POLLS   75%: Take Country Back From Rich &amp; Powerful https://t.co/nIBXu9aHl4  #ElectionNight https://t.
allisg|WinterAntiques|0.3612|0.0|0.872|0.128|"RT @WinterAntiques: The chicest accessory on Election Day? An ""I voted"" sticker.  #ElectionDay #Election2016 #portrait  Courtesy of Ro"
mezthlyy|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
EscapeWithTessa|twitter|0.0|0.0|1.0|0.0|This election reminds me of https://t.co/Wj8aXbYxXL
lafrogh|TheEconomist|0.0|0.0|1.0|0.0|RT @TheEconomist: Alaska's native Americans are traditionally under-represented in elections https://t.co/VjvDTwpXk3
lafrogh|economist|0.0|0.0|1.0|0.0|RT @TheEconomist: Alaska's native Americans are traditionally under-represented in elections https://t.co/VjvDTwpXk3
Manda_Guards|LoveYourMelon|0.6239|0.0|0.823|0.177|RT @LoveYourMelon: Beanies + Ballots = A Successful Election DayCheck out our new products as you wait in line to cast your ballot!https:
allenvollbrecht|wikileaks|-0.5994|0.178|0.822|0.0|RT @wikileaks: US presidential candidate @DrJillStein (Greens) draws attention to Obama's war on whistleblowers in election eve PR https://
allenvollbrecht||-0.5994|0.178|0.822|0.0|RT @wikileaks: US presidential candidate @DrJillStein (Greens) draws attention to Obama's war on whistleblowers in election eve PR https://
Benross75|Benross75|0.6239|0.0|0.806|0.194|"RT @Benross75: .@BretBaier @realDonaldTrump  Trump is up in Florida and North Carolina, let's win this election Tomorrow People!"
Akexfromtarget|MikeDrucker|0.0|0.0|1.0|0.0|RT @MikeDrucker: Yo can we have a big smash bros tournament on your screens after the election https://t.co/Zda4wZIh88
Akexfromtarget|twitter|0.0|0.0|1.0|0.0|RT @MikeDrucker: Yo can we have a big smash bros tournament on your screens after the election https://t.co/Zda4wZIh88
jojo_cha_1|greta|0.6369|0.0|0.84|0.16|"RT @greta: Would love to see some anchoring of election coverage from mid west/west USA..would remind people this is a big country, not jus"
amezalim|BernieSanders|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
amezalim|twitter|0.4404|0.0|0.847|0.153|RT @BernieSanders: Today is an election of enormous consequence. I hope everybody gets out to vote. #ElectionDay https://t.co/JYYunxLO2R
GCC_legal|reuters|0.0|0.0|1.0|0.0|RT ReutersPolitics: Former President George W. Bush does not cast vote for president https://t.co/GvFhbiQ1uc
bgordian01|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
mvjennings|wlunews|0.4926|0.0|0.738|0.262|@wlunews Fond memories of producing Channel 9 election coverage in 1992!
oldwalren|LaurenJauregui|0.6892|0.0|0.738|0.262|RT @LaurenJauregui: Freakin out about Election Day lol make sure you all go out and VOTEEEEE TOMORROW!! #imwithHER
_TheMayor|Bencjacobs|0.0|0.0|1.0|0.0|RT @Bencjacobs: Cash bar at trump election night event
loriwitherell|greggutfeld|0.0|0.0|1.0|0.0|RT @greggutfeld: my monologue on how to react to the election: https://t.co/y4DgRFkbpj
loriwitherell|video|0.0|0.0|1.0|0.0|RT @greggutfeld: my monologue on how to react to the election: https://t.co/y4DgRFkbpj
Vianney678|CNN|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
Vianney678|twitter|0.0|0.0|1.0|0.0|RT @CNN: Stand by for #CNNElection projectionhttps://t.co/15RGLqdxpK#ElectionNight https://t.co/Ty5O1defYU
ButeraFtDinah|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
ButeraFtDinah|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
mehdifoundation|medium|0.0|0.0|1.0|0.0|#Terrorism and the Presidential Election: https://t.co/f3gu5ZIsCM #HillaryClinton #DonaldTrump #ImWithHer #ElectionNight #USA
mrbobfan11|twitter|0.0|0.0|1.0|0.0|Watching the #election https://t.co/SMHtaXqlU3
isaganimeliton|wsj|0.0|0.0|1.0|0.0|Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/WR2biShRT3  #Election2016... https://t.co/wPUSlPrk1M
alxdark|GoAngelo|0.0|0.0|1.0|0.0|"RT @GoAngelo: Election Night 2012Actual ResultsObama: 65,915,795Romney: 60,933,504 https://t.co/dtD8WwpAd6"
alxdark|twitter|0.0|0.0|1.0|0.0|"RT @GoAngelo: Election Night 2012Actual ResultsObama: 65,915,795Romney: 60,933,504 https://t.co/dtD8WwpAd6"
scott_isler|CNNPolitics|0.0|0.0|1.0|0.0|Election 2016: Live coverage @CNNPolitics https://t.co/R6BBTXeGj8
scott_isler|cnn|0.0|0.0|1.0|0.0|Election 2016: Live coverage @CNNPolitics https://t.co/R6BBTXeGj8
AdamHasner|LRSpies|0.304|0.079|0.757|0.164|RT @LRSpies: @katiepack @Timodc please tweet often so I don't have to bother @cspiesdc He ignores me &amp; just sends me this link https://t.c
AdamHasner||0.304|0.079|0.757|0.164|RT @LRSpies: @katiepack @Timodc please tweet often so I don't have to bother @cspiesdc He ignores me &amp; just sends me this link https://t.c
wptweetmachine|tricks4|0.4019|0.0|0.816|0.184|The kitten mindfulness video you need to help you keep your electionchill https://t.co/ZhRZjXnKrw
election_votes|Hxrnet|0.0772|0.0|0.894|0.106|RT @Hxrnet: I want to see who you guys are favoring/voting for.. Pick.
NouveauGlass|fivethirtyeight|0.2023|0.0|0.899|0.101|How important is Florida? (Polls in the eastern part of the stateclose in a few minutes.) If https://t.co/sV5z9s1Pu9
legumehs|CherOfficiaI|0.6633|0.0|0.783|0.217|RT @CherOfficiaI: IF TRUMP WINS THE ELECTION   I AM MOVIN OUT OF THE COUNTRY  GOODBYE AMERICA HELLO  CALIFORNIA
friwaysblog|haaretzcom|0.7096|0.0|0.772|0.228|RT @haaretzcom: Polls in parts of Florida are about to close. Will the Muslim vote help hand Florida to Clinton? https://t.co/oqUgaoUu5I ht
friwaysblog|haaretz|0.7096|0.0|0.772|0.228|RT @haaretzcom: Polls in parts of Florida are about to close. Will the Muslim vote help hand Florida to Clinton? https://t.co/oqUgaoUu5I ht
leahh617|PatrickRothfuss|0.0|0.0|1.0|0.0|RT @PatrickRothfuss: Reminder: In Wisconsin you can register to vote at your polling place on election day.For real. Same-day registratio
dinobuttz|lizacsg|0.0|0.0|1.0|0.0|"RT @lizacsg: sometimes the election gets me down. but then, cheese. https://t.co/HG8AFl3igl"
dinobuttz|twitter|0.0|0.0|1.0|0.0|"RT @lizacsg: sometimes the election gets me down. but then, cheese. https://t.co/HG8AFl3igl"
TAKEBACKOCH|miamiherald|0.0|0.0|1.0|0.0|RT: Shooting in California leaves two polling places on lock down https://t.co/0gTB1hAXzz https://t.co/u6h0xMRf8A via MiamiHerald
LokoAzzE_man|twitter|0.0|0.0|1.0|0.0|Ya WCW thought inauguration and Election Day was the same day https://t.co/mJJBb5fFYe
Mom74548299|roycan79|0.0|0.0|1.0|0.0|"RT @roycan79: UPDATE: Election will in all probability go down to the WIRE, so we NEED EVERY LAST VOTE for #TRUMP!  PUSH YOURSELF! GO VOTE!"
marshray|NPR|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
marshray|npr|0.4019|0.0|0.863|0.137|RT @NPR: Los Angeles authorities say two polling locations are closed due to an active shooter situation. https://t.co/C7Y1uiDgpf
delawareonline|delawareonline|0.0|0.0|1.0|0.0|#ElectionNight is finally here: What you need to know now. https://t.co/0PiKJA9qXI #voteDE
bigbrownie167|NounouBby|0.8068|0.0|0.751|0.249|RT @NounouBby: I mean the election may be over tonight but I'll never forget how racist some of y'all are so are you really safe????
domedog311|"Always_Trump,#TrumpArmy,"|-0.4101|0.155|0.845|0.0|"@Always_Trump,#TrumpArmy, #TrumpTrain, @BigStick2013,@ChrisCoon4 I've never been so nervous waiting for election night returns. Much on line"
MikeDarnay|HockeyBabbler|0.2748|0.0|0.905|0.095|"RT @HockeyBabbler: There will almost certainly be people who stay at home because of this, and that can sway an election."
sabrobidoux|ABC|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
sabrobidoux|abcnews|-0.0258|0.096|0.812|0.092|RT @ABC: Scores of people wait in line to say thank you at the grave of voting rights activist Susan B. Anthony. https://t.co/IKTN8J2oeN ht
thattattedupguy|riverandmal|-0.5423|0.241|0.759|0.0|@riverandmal This would be a real bad election for them to elected anyone.
obeyyurTHURST|PresidentJalen|-0.4939|0.39|0.61|0.0|RT @PresidentJalen: Election Night Lowkey scary
ConnieInAmerica|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
ConnieInAmerica|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Election Day is almost over. Dont waitgo vote now! Confirm where you vote at https://t.co/jfd3CXLD1s https://t.co/Iv
myia_rae|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
myia_rae|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
silverfoxmedia1|FredZeppelin12|0.25|0.0|0.895|0.105|RT @FredZeppelin12: DRUDGE: ELECTION WILL BE DECIDED BY EVENING VOTERS. Advantage #Trump. Evening voters are evening voters because t
politicallynate|NateSilver538|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
politicallynate|fivethirtyeight|0.4767|0.121|0.603|0.276|"RT @NateSilver538: If Clinton wins Florida, her chances will shoot up to about 93%. https://t.co/ZUCgeSJ5eP"
loneevolution|Princessofwifi|-0.5574|0.295|0.705|0.0|RT @Princessofwifi: Forget the US election the Uk is facing a bigger problem  https://t.co/PErV4k692k
loneevolution|twitter|-0.5574|0.295|0.705|0.0|RT @Princessofwifi: Forget the US election the Uk is facing a bigger problem  https://t.co/PErV4k692k
andrewkmorse|CNET|0.0|0.0|1.0|0.0|Can social media call the election? https://t.co/mh9iX9EXCD via @CNET #Election2016 #ElectionNight
andrewkmorse|cnet|0.0|0.0|1.0|0.0|Can social media call the election? https://t.co/mh9iX9EXCD via @CNET #Election2016 #ElectionNight
TheMusicMamaB|Debramax|0.0|0.0|1.0|0.0|"RT @Debramax: BREAKING : African American Female Trump Exec Says ""Blacks Will Swing the Election to Trump"" https://t.co/ZvNWKBhDeE"
TheMusicMamaB|truthfeed|0.0|0.0|1.0|0.0|"RT @Debramax: BREAKING : African American Female Trump Exec Says ""Blacks Will Swing the Election to Trump"" https://t.co/ZvNWKBhDeE"
JohnProchello|LifeAsRednecks|0.0|0.0|1.0|0.0|RT @LifeAsRednecks: Election Prediction: Democrats take an early lead until Republicans finally get off work to go and vote
gabipjunkes|Telegraph|-0.6486|0.223|0.777|0.0|RT @Telegraph: #ElectionNight One person is reportedly dead after a shooting in California near a polling station https://t.co/CJCBsKKKNE
gabipjunkes|telegraph|-0.6486|0.223|0.777|0.0|RT @Telegraph: #ElectionNight One person is reportedly dead after a shooting in California near a polling station https://t.co/CJCBsKKKNE
princess_nanas|picudoooooo|-0.6597|0.355|0.645|0.0|"RT @picudoooooo: After the election, we're fucked either way"
LGarchomp|Crunchyroll|-0.2244|0.12|0.793|0.087|"RT @Crunchyroll: Today's ELECTION DAY in the US, make sure to vote!...but if you're tired of 538 electoral maps, we have one that's a"
WhosGoneGalt|An0nRav|-0.7351|0.341|0.659|0.0|RT @An0nRav: Report fraud or disruptions at polling locationsVoter Assistance Hotline:at (844) 332-2016Or online:https://t.co/xbhHANrIB
WhosGoneGalt|t|-0.7351|0.341|0.659|0.0|RT @An0nRav: Report fraud or disruptions at polling locationsVoter Assistance Hotline:at (844) 332-2016Or online:https://t.co/xbhHANrIB
MartinCartermc3|JamesOKeefeIII|0.7027|0.0|0.779|0.221|"RT @JamesOKeefeIII: WOW! Caught more #VoterFraud in N Philly. Election workers caught BREAKING THE LAW. #VeritasIsEverywhere Stay tuned, co"
Chulaa54|2inchesOfDoom|-0.5574|0.286|0.714|0.0|RT @2inchesOfDoom: I can't wait till this election shit over with.
BillyH_mdr|Venice311|0.0772|0.0|0.933|0.067|"RT @Venice311: If you want the realtime results for the LA County Election stuff + POTUS NEVAUX, clicky clicky: https://t.co/gOA4S7cRos"
BillyH_mdr|lavote|0.0772|0.0|0.933|0.067|"RT @Venice311: If you want the realtime results for the LA County Election stuff + POTUS NEVAUX, clicky clicky: https://t.co/gOA4S7cRos"
Go_gedem|ABC|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
Go_gedem|t|-0.4404|0.121|0.879|0.0|"RT @ABC: Trump, Clinton are both in Midtown Manhattan tonight, watching the results come in just a block away from each other https://t.co/"
HectorPooley|linkis|0.802|0.0|0.613|0.387|"Reuters/Ipsos Exit Poll: 3 in 4 Think Economy 'Rigged' for 'Rich and Powerful,' Want 'Strong Leader' - Breitbart https://t.co/eboeh1fExx"
BrickStOxford|twitter|0.508|0.0|0.785|0.215|Watch the election unfold right here! Special edition red or blue trashcans! https://t.co/ULhy481iNW
DrDrizzleh|wolfieraps|0.7865|0.0|0.783|0.217|RT @wolfieraps: If trump wins the election today who wants to come back to Canada with me? LIKE this tweet so I know to buy you an airplane
wxgarrett|ActionNewsJax|0.4019|0.0|0.838|0.162|RT @ActionNewsJax: NOW: Watch our special election coverage on FOX30 or Facebook Live: https://t.co/WqUi3oMIUg https://t.co/lscZNdoOuh
wxgarrett|facebook|0.4019|0.0|0.838|0.162|RT @ActionNewsJax: NOW: Watch our special election coverage on FOX30 or Facebook Live: https://t.co/WqUi3oMIUg https://t.co/lscZNdoOuh
BellaBootySDMN|memetribute|-0.6371|0.259|0.741|0.0|RT @memetribute: LEAKED RESULTS OF TONIGHTS ELECTION IN WHICH JEB FIXED IT!!!! https://t.co/dRJafaQaQU
BellaBootySDMN|twitter|-0.6371|0.259|0.741|0.0|RT @memetribute: LEAKED RESULTS OF TONIGHTS ELECTION IN WHICH JEB FIXED IT!!!! https://t.co/dRJafaQaQU
alehra_|carwash54|0.7085|0.0|0.734|0.266|"RT @carwash54: Me @ the beginning of the election: Ain't no way America letting a cheeto become president. lol what a joke Me November 7,"
nicky02345|washingtonpost|-0.3818|0.167|0.833|0.0|Jon Stewart joins Stephen Colbert to slam Trump once more on election eve https://t.co/7LNghckdi9
zatheteacher|mashable|0.0|0.0|1.0|0.0|America gets lit: The Lite Brite guide to election results https://t.co/dSsH54haDn
CheetahPizzas|OPB|-0.3818|0.148|0.852|0.0|"RT @OPB: At Susan B. Anthony's Grave, visiting hours extended for election day crowds  https://t.co/KWJS1XealL https://t.co/YItRaU3xO1"
CheetahPizzas|opb|-0.3818|0.148|0.852|0.0|"RT @OPB: At Susan B. Anthony's Grave, visiting hours extended for election day crowds  https://t.co/KWJS1XealL https://t.co/YItRaU3xO1"
_GBR2|GovMikeHuckabee|0.4019|0.0|0.844|0.156|"RT @GovMikeHuckabee: Analysts say election will be determined by after-work voters. If you have a job, or ever want one, go vote Trump."
HareshShah2014|clusterstock|0.5719|0.0|0.821|0.179|RT @clusterstock: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/x7Sl4pgVPC https://t.co/Q
HareshShah2014|businessinsider|0.5719|0.0|0.821|0.179|RT @clusterstock: WORLD'S BIGGEST HEDGE FUND: Stock markets around the world will tank if Trump wins https://t.co/x7Sl4pgVPC https://t.co/Q
iamprikle|asunnydisposish|-0.2263|0.076|0.924|0.0|"RT @asunnydisposish: As someone who can't vote today but will still be affected by the election results, I urge you to not throw away your"
Gungledink|democracynow|0.0|0.0|1.0|0.0|WATCH: Election Night 2016 Coverage with Democracy Now! https://t.co/Jr2wo02BrE via @democracynow
Gungledink|democracynow|0.0|0.0|1.0|0.0|WATCH: Election Night 2016 Coverage with Democracy Now! https://t.co/Jr2wo02BrE via @democracynow
CalebBrankle|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
k8linsucks|repjohnlewis|0.0|0.0|1.0|0.0|"RT @repjohnlewis: Do not give up, give in, or give out. You must do what it takes to make your voice heard and cast your ballot in this ele"
Aljaberzoon|nytimes|0.0|0.0|1.0|0.0|RT @nytimes: Who will you vote for? Get the facts on the NYTimes Election Guide. https://t.co/rByycsGXxI
Aljaberzoon|itunes|0.0|0.0|1.0|0.0|RT @nytimes: Who will you vote for? Get the facts on the NYTimes Election Guide. https://t.co/rByycsGXxI
MrKline_EdTech|mrhushistory|-0.2377|0.093|0.907|0.0|"RT @mrhushistory: @TecumsehJrHigh students I'll be your source (and way more fun!!) for unbiased Election 2016 coverage, news &amp; insights.Go"
SzulimJula|RachelAndJun|-0.3384|0.23|0.77|0.0|RT @RachelAndJun: So nervous about the election I can't sleep
sheilajsampson|JamesOKeefeIII|-0.5423|0.132|0.868|0.0|"RT @JamesOKeefeIII: We just caught election officials telling people who to vote for, crime Under 25 PS 3031.11. I will tag both you and @D"
paulrlanni|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
JoshGellers|WJCTJax|0.0|0.0|1.0|0.0|Prepping for live #election coverage @WJCTJax w/ @MelissainJax! #ElectionNight @NPR https://t.co/JSIhFhYcY4
JoshGellers|twitter|0.0|0.0|1.0|0.0|Prepping for live #election coverage @WJCTJax w/ @MelissainJax! #ElectionNight @NPR https://t.co/JSIhFhYcY4
Rosenchild|CNNPolitics|0.0|0.0|1.0|0.0|RT @CNNPolitics: Women in pantsuits send a message on #ElectionDay https://t.co/s2GZLEg889 https://t.co/RphWoVplBU
Rosenchild|cnn|0.0|0.0|1.0|0.0|RT @CNNPolitics: Women in pantsuits send a message on #ElectionDay https://t.co/s2GZLEg889 https://t.co/RphWoVplBU
SaharaTV1|lizgrossman87|0.0|0.0|1.0|0.0|RT @lizgrossman87: Check out @SaharaTV1's #uselection coverage of the election @haingovalencia https://t.co/POaV1ynOrq. #Nov8AfricanEdition
SaharaTV1|youtube|0.0|0.0|1.0|0.0|RT @lizgrossman87: Check out @SaharaTV1's #uselection coverage of the election @haingovalencia https://t.co/POaV1ynOrq. #Nov8AfricanEdition
peejaybee|daveweigel|0.1027|0.118|0.746|0.136|"RT @daveweigel: With less than 1% of my post-election diet underway, I can confidently report that I will lose 50 pounds."
cheycll|conserv_tribune|0.0|0.0|1.0|0.0|RT @conserv_tribune: BREAKING: All Election Systems Are Down in Swing State of Colorado https://t.co/xCpH7pZEkY #tcot https://t.co/JNZLA8
cheycll|conservativetribune|0.0|0.0|1.0|0.0|RT @conserv_tribune: BREAKING: All Election Systems Are Down in Swing State of Colorado https://t.co/xCpH7pZEkY #tcot https://t.co/JNZLA8
SnoVitKatt|djajiprime|0.5267|0.0|0.779|0.221|"RT @djajiprime: Enjoying the election coverage with #TYTlive, you can watch too:https://t.co/TwdOpIsuaj#ElectionNight https://t.co/l6cllx"
SnoVitKatt|youtube|0.5267|0.0|0.779|0.221|"RT @djajiprime: Enjoying the election coverage with #TYTlive, you can watch too:https://t.co/TwdOpIsuaj#ElectionNight https://t.co/l6cllx"
ambree_cuyler|quote_friends|0.3612|0.0|0.706|0.294|RT @quote_friends: election got me like https://t.co/ZuZ8kMVSJM
ambree_cuyler|twitter|0.3612|0.0|0.706|0.294|RT @quote_friends: election got me like https://t.co/ZuZ8kMVSJM
HANN_itToAh|chungaah|0.3818|0.122|0.667|0.211|RT @chungaah: Not even worried about the election Ik who gonna win Hillary obviously 
ardie2pt0|BernieSanders|0.6705|0.0|0.776|0.224|RT @BernieSanders: I can't fill in for every worker today. Election Day should be a national holiday so that everyone has the opportunity t
PTicks|WSJ|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
PTicks|wsj|0.0|0.0|1.0|0.0|RT @WSJ: Polls close in six states at 7 p.m. EST. Follow along for live updates: https://t.co/reNrPgubQ6  #Election2016 https://t.co/pz4iZ
Mom_Im_Sorry|jeffpeartshow|0.0|0.0|1.0|0.0|"RT @jeffpeartshow: EP: 45 A VOTE FOR CHANGE We finally let Gary talk about the election + a $5,000 Cheeto.https://t.co/sDgvK84HSf#Podern"
outsidethewire2|mikeroman|0.0|0.0|1.0|0.0|"RT @mikeroman: Hearing in Philly: Pollwatcher testifying that Election Judge ""pushed"" him out of the poling place."
AmIThatBad|UpshotNYT|0.5859|0.0|0.725|0.275|RT @UpshotNYT: When will we know we have a winner? https://t.co/1pMJXK7mS4 https://t.co/B87hwbBQZy
AmIThatBad|nytimes|0.5859|0.0|0.725|0.275|RT @UpshotNYT: When will we know we have a winner? https://t.co/1pMJXK7mS4 https://t.co/B87hwbBQZy
young_maymay|HuffPostPol|0.0|0.0|1.0|0.0|RT @HuffPostPol: And follow our live analysis right here: https://t.co/PmkRCmLxFx #election https://t.co/7CSTTdsvCp
young_maymay|huffingtonpost|0.0|0.0|1.0|0.0|RT @HuffPostPol: And follow our live analysis right here: https://t.co/PmkRCmLxFx #election https://t.co/7CSTTdsvCp
CxntBe_Tamed|bxddaddiction|0.7184|0.0|0.75|0.25|RT @bxddaddiction: Come to the election party tonight at OT doors open at 8 free shot of ciroc for voters https://t.co/ZmmZqcKVZ9
CxntBe_Tamed|twitter|0.7184|0.0|0.75|0.25|RT @bxddaddiction: Come to the election party tonight at OT doors open at 8 free shot of ciroc for voters https://t.co/ZmmZqcKVZ9
TheRogueelement|realDonaldTrump|0.2124|0.0|0.931|0.069|"RT @realDonaldTrump: Don't let up, keep getting out to vote - this election is FAR FROM OVER! We are doing well but there is much time left"
SquidlyM|memeprovider|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
SquidlyM|twitter|0.0|0.0|1.0|0.0|RT @memeprovider: got my election sticker https://t.co/EBknYdpVzU
charlotteole1|denverpost|0.0|0.0|1.0|0.0|"RT @denverpost: LIVE BLOG: Live #Election2016 updates, results, stories, and full #copolitics coverage from across Colorado https://t.co/SJ"
charlotteole1|t|0.0|0.0|1.0|0.0|"RT @denverpost: LIVE BLOG: Live #Election2016 updates, results, stories, and full #copolitics coverage from across Colorado https://t.co/SJ"
livenewscloud|livenewscloud|0.296|0.0|0.885|0.115|#BREAKING Watch live: Join @livenewscloud during historic election as first results come in in 2mins LIVESTREAM &gt;&gt;&gt; https://t.co/ZWqnCp3cek
livenewscloud|livenewschat|0.296|0.0|0.885|0.115|#BREAKING Watch live: Join @livenewscloud during historic election as first results come in in 2mins LIVESTREAM &gt;&gt;&gt; https://t.co/ZWqnCp3cek
