User|Original_User/Web|Compound|Negative|Neutral|Positive|Tweet
_bigpharma|RicheyCollazo|0.8356|0.0|0.603|0.397|RT @RicheyCollazo: white women: Hillary Clintons win is a win for women!me: WHICH WOMEN?  https://t.co/FONDX957Gy
_bigpharma|twitter|0.8356|0.0|0.603|0.397|RT @RicheyCollazo: white women: Hillary Clintons win is a win for women!me: WHICH WOMEN?  https://t.co/FONDX957Gy
br1xanna|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
gelegwen|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
gelegwen|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
Larkell_|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
fredbauerblog|nationalreview|0.0|0.0|1.0|0.0|"Before the deluge of results, I'll reiterate this: Our republic will survive whatever the result. https://t.co/TUW7beveWb"
RespectOurFlag2|WDFx2EU8|-0.6739|0.232|0.768|0.0|RT @WDFx2EU8: WIDESPREAD VOTER FRAUD: Philadelphia Democrats Pass Out Pro-Hillary Brochures At Polling Sites (VIDEO) https://t.co/7w2LzjPIYc
RespectOurFlag2|americanlookout|-0.6739|0.232|0.768|0.0|RT @WDFx2EU8: WIDESPREAD VOTER FRAUD: Philadelphia Democrats Pass Out Pro-Hillary Brochures At Polling Sites (VIDEO) https://t.co/7w2LzjPIYc
suleikamenaa|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
suleikamenaa|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Tiph_Seven|parksandrecnbc|0.0|0.0|1.0|0.0|"Hillary got to come out to ""Get on your feet"" one time for @parksandrecnbc #ClintonKnope"
sherrymisner|dawg_lb|0.0|0.0|1.0|0.0|"RT @dawg_lb: Hillary R Clinton,YOU SHOULD NEVER BE ABLE TO LOOK AT YOURSELF IN THE MIRROR!!!!!!!VOTE AS FAST AS YOU CAN!!!!!!!!!!TRUM"
Isaiah1337|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
parettijacob|REALBrianStreng|0.7096|0.0|0.789|0.211|RT @REALBrianStreng: Joke is on Hillary if she wins the election because that means she has to sit at the desk Monica was under
nicholas51|newsmax|0.0|0.0|1.0|0.0|"RT @newsmax: With 1% of the vote in for Kentucky, Trump is holding a steady lead over Hillary Clinton. #ElectionNight #myvote2016 https://t"
nicholas51||0.0|0.0|1.0|0.0|"RT @newsmax: With 1% of the vote in for Kentucky, Trump is holding a steady lead over Hillary Clinton. #ElectionNight #myvote2016 https://t"
shelbghughes|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
shelbghughes|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
_SAVE_AMERICA|WayneDupreeShow|-0.296|0.136|0.864|0.0|RT @WayneDupreeShow:  Huckabee: Hillary Has No Empathy For The Working Class https://t.co/NEEjhHx6Zy #DrainTheSwamp #TrumpTrain https://t.
_SAVE_AMERICA|newsninja2012|-0.296|0.136|0.864|0.0|RT @WayneDupreeShow:  Huckabee: Hillary Has No Empathy For The Working Class https://t.co/NEEjhHx6Zy #DrainTheSwamp #TrumpTrain https://t.
feltonewt|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
blurrygambino|twitter|0.128|0.169|0.635|0.196|When you realize that we're screwed if trump or Hillary wins the election https://t.co/5ULRBFJVIR
andBridget|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
blujayva|JudicialWatch|0.2023|0.0|0.909|0.091|RT @JudicialWatch: Hillary and many of her top aides treated the court process with contempt.View our Weekly Update here.https://t.co/qjW
courtalexandra_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
itssallymarie|AfroGumOfficiaI|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
itssallymarie|twitter|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
_Kareem12|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
yanesque|sassytbh|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
yanesque|twitter|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
4peaks94|mitchellvii|-0.7645|0.32|0.68|0.0|"RT @mitchellvii: Based upon exits, voters very unhappy with big money corruption.  That's bad for Hillary."
DrThomasPaul|DrThomasPaul|-0.1531|0.164|0.701|0.136|"RT @DrThomasPaul: .@HillarysAmerica is one of division, crime, #pharma &amp; riots.It's good for corrupt #BigBusiness.#gmo #Hillary #Trumphttp"
_KFrye|EvanFoerster|0.3612|0.0|0.615|0.385|RT @EvanFoerster: @_KFrye u like hillary?
erekaarmstead|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
erekaarmstead|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
thiboteirlinck|DaiIyRap|0.0772|0.0|0.86|0.14|RT @DaiIyRap: Hillary Clinton doing the Mannequin Challenge https://t.co/yZXFZ1hNrn
thiboteirlinck|twitter|0.0772|0.0|0.86|0.14|RT @DaiIyRap: Hillary Clinton doing the Mannequin Challenge https://t.co/yZXFZ1hNrn
BeatsBy777|UglyGod|-0.5106|0.121|0.879|0.0|RT @UglyGod: It means yall shoulda fuckin listened &amp; kept Bernie Sanders as an option cause now we all look dumb af choosing between Hillar
HeelStCloud|Rokkaaaaa|-0.6705|0.287|0.599|0.114|"RT @Rokkaaaaa: I laugh at people whose main beef with Hillary is lying. Dude people lie everyday. Today, I lied and blamed metro for being"
LeighaCrumpler|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
LeighaCrumpler|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
TarnTawanxx|billboard|0.0|0.0|1.0|0.0|RT @billboard: Mother Monster wants you to vote.   https://t.co/988SkvrQOx https://t.co/CHliI37Ymk
TarnTawanxx|billboard|0.0|0.0|1.0|0.0|RT @billboard: Mother Monster wants you to vote.   https://t.co/988SkvrQOx https://t.co/CHliI37Ymk
ruthe_susan|Wil_Johnson1|0.0|0.0|1.0|0.0|"RT @Wil_Johnson1: In Kentucky and Indiana with just a little over 3% reporting, Trump is getting 2-1 votes over Hillary https://t.co/4wCD0Q"
ruthe_susan|t|0.0|0.0|1.0|0.0|"RT @Wil_Johnson1: In Kentucky and Indiana with just a little over 3% reporting, Trump is getting 2-1 votes over Hillary https://t.co/4wCD0Q"
JenTromans|Alex_Hxrrison|0.3291|0.0|0.895|0.105|"RT @Alex_Hxrrison: If Hillary wins then she is the first F president. Oops should've been female but the ""emale"" got deleted #ElectionDay #"
atf13atf|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
keluttcu|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
czareah_|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
czareah_|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
dgraz007|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
dgraz007|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
sunshinejilly45|YoungDems4Trump|-0.0258|0.14|0.725|0.135|RT @YoungDems4Trump: Hillary should be tried for Treason. Not run for the President of the United States.#ElectionDay#MyVote2016
MarioHazelwood|ZachAJacobson|0.8625|0.0|0.676|0.324|"RT @ZachAJacobson: Yes, I voted Hillary. You voted Trump? Nice. Won't change how I, or anybody else should view you. Great thing about Amer"
coolstuffbynawk|philsadelphia|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
coolstuffbynawk|twitter|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
LESTERHICKEYS|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
LESTERHICKEYS|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
ninabautista|AFP|0.0|0.0|1.0|0.0|"RT @AFP: A large Hillary for America sign is displayed at the Jacob K. Javits Center in New York, where Clinton's #ElectionNight event is h"
carybaskin|2ALAW|-0.4404|0.231|0.602|0.167|"RT @2ALAW: It's truly a sad day in America when we dismiss all the corruption, voting fraud committed as ""just politics""#Hillary is disqu"
CDavidlynn|lifenews|0.8074|0.0|0.52|0.48|Hillary Clinton: I Want a Supreme Court Justice Who Will Uphold Unlimited Abortion https://t.co/UfgCOjWXzC
AMGR84|claireholt|0.0|0.0|1.0|0.0|@claireholt @elenaahh20 I VOTED FOR HILLARY!! I'AM WITH HER! VOTE GUYS!
kielymarie26|misheardhamilto|0.0|0.0|1.0|0.0|RT @misheardhamilto: and if you were to ask me who i'd promote?hillary has my vote #ElectionDay
Kahless_72|gerfingerpoken|-0.5106|0.202|0.798|0.0|RT @gerfingerpoken: Hillary Clinton's Failing Health a Real Concern https://t.co/OkDpwx6Jgf - #PJNET 999 - American Thinker - https://t.co/
Kahless_72|americanthinker|-0.5106|0.202|0.798|0.0|RT @gerfingerpoken: Hillary Clinton's Failing Health a Real Concern https://t.co/OkDpwx6Jgf - #PJNET 999 - American Thinker - https://t.co/
semperadlucum|cnn|-0.0018|0.108|0.784|0.108|"@cnn Dont worry u media made it very clear who u wanted as POTUS. Hillary is ur baby and u wanted to,protect her all the way."
KeepEmAccntable|weknowwhatsbest|0.8225|0.0|0.688|0.312|"RT @weknowwhatsbest: I wish Hillary's ""Our Kids Are Watching"" speech would have been followed by a lovely song from her #1 supporter Jay Z."
zuvysypemufyw|itegistry|0.5859|0.0|0.703|0.297|Hillary - https://t.co/J433FXzTyd Stock Market Is Leaning Toward a Hillary Clinton Win
natkovacevich|LifeAsRednecks|0.6124|0.0|0.773|0.227|RT @LifeAsRednecks: Votin for Hillary just because shes a woman is like drinkin antifreeze just because it looks like Gatorade.
jimmybelshe|DRUDGE_REPORT|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
jimmybelshe|businessinsider|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
bear_oyo|ProfessorF|0.8225|0.0|0.703|0.297|"RT @ProfessorF: Wow another example of Hillary's ""superior"" ground game. That's brilliant. Having election officials tell people who to vot"
gruvvywave|c0nvey|0.0|0.0|1.0|0.0|Hillary Clinton is privately against gay marriage https://t.co/vgWFzoErKT by #wikileaks via @c0nvey
gruvvywave|linkis|0.0|0.0|1.0|0.0|Hillary Clinton is privately against gay marriage https://t.co/vgWFzoErKT by #wikileaks via @c0nvey
LenahanChris|weknowwhatsbest|-0.3804|0.166|0.834|0.0|RT @weknowwhatsbest: Exit polling shows that Hillary has completely lost the 3rd trimester vote.
iamronaldpaul|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @Slate @votecastr @LilSteelerGirl @DebAlwaystrump @Kerri1111 TRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLID
ecwpunk81|HillaryforOH|0.0|0.0|1.0|0.0|RT @HillaryforOH: Ohio polls are open until 7:30pmfind your voting location at https://t.co/2otkpVPJlw and go cast your ballot for Hillary
ecwpunk81|iwillvote|0.0|0.0|1.0|0.0|RT @HillaryforOH: Ohio polls are open until 7:30pmfind your voting location at https://t.co/2otkpVPJlw and go cast your ballot for Hillary
chrgdup1973|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
iDreamRihanna|MTVstyle|0.0|0.0|1.0|0.0|RT @MTVstyle: Rihanna wore a t-shirt of HERSELF wearing a Hillary Clinton t-shirt because SHE IS THE STYLE ICON OUR NATION NEEDS:https://
iDreamRihanna||0.0|0.0|1.0|0.0|RT @MTVstyle: Rihanna wore a t-shirt of HERSELF wearing a Hillary Clinton t-shirt because SHE IS THE STYLE ICON OUR NATION NEEDS:https://
allycook108|laneonme|0.7964|0.0|0.755|0.245|RT @laneonme: and if you vote hillary make sure you tell all your friends and family in the military that you support her &amp; what she did wi
patrickjalbino|JoyAnnReid|0.3182|0.0|0.887|0.113|RT @JoyAnnReid: Hillary Clinton being tied among white voters with a college degree is actually a huge swing toward Democrats. #ExitPolls
GJoelChury|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
BustosBella|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
hostagehoosier|mamaswati|-0.3182|0.103|0.897|0.0|@mamaswati lady with the hillary sticker looked genuinely shocked when i glared at her after she asked if I wanted a sample dem ballot.
_3Digital|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_3Digital|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
princessle4h|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
princessle4h|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
AmbieeJojo|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
AmbieeJojo|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Lenka_|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
jezzybees|ashiebaker|-0.4574|0.136|0.864|0.0|"Chris Wallace just asked ""what if Hillary flips GA?""  @ashiebaker and @MelaninDSass will lose their chill is what will happen!"
sbca80|TheEconomist|-0.7506|0.39|0.61|0.0|RT @TheEconomist: Donald Trump's reckless foreign policy could unleash chaos https://t.co/kJPHr47hHn https://t.co/VhOjRhE6br
sbca80|economist|-0.7506|0.39|0.61|0.0|RT @TheEconomist: Donald Trump's reckless foreign policy could unleash chaos https://t.co/kJPHr47hHn https://t.co/VhOjRhE6br
llylahh__|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
llylahh__|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
FranCarmichael|NathanZed|0.5267|0.0|0.848|0.152|RT @NathanZed: my 7 year old cousin just now: is Hellen Keller winning me: whatcousin: Hellen Kellerme: Hillary Clinton? cousin: I dont
_ariannneeezy|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
_ariannneeezy|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
HansonbooRiah|jozenc|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
HansonbooRiah|twitter|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
_KrissyGomez|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Bungalow0|anonymous585446|0.0|0.0|1.0|0.0|@anonymous585446 Guam. Hillary 72%
DriggersJudy|suziedaud|0.0|0.0|1.0|0.0|"RT @suziedaud: #DNCLeak2 Hillary's staffers discussing Bill &amp; Epsteins #LolitaExpress with underage girls on way to ""Orgy Island""https://"
DriggersJudy||0.0|0.0|1.0|0.0|"RT @suziedaud: #DNCLeak2 Hillary's staffers discussing Bill &amp; Epsteins #LolitaExpress with underage girls on way to ""Orgy Island""https://"
iridescentnoir|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
iridescentnoir|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
russmove|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
twinkIouis|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
twinkIouis|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
TheMadHessian|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
TheMadHessian|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Thompson1226||0.0|0.0|1.0|0.0|"I voted for Hillary, don't @ me"
annyglop23|Latina_pe|0.0|0.0|1.0|0.0|RT @Latina_pe: Boca de urna- New Hampshire: Donald Trump: 52% Hillary Clinton: 41% #EleccionesEEUU #ElectionDay https://t.co/uhnyqN3ZuC
annyglop23|twitter|0.0|0.0|1.0|0.0|RT @Latina_pe: Boca de urna- New Hampshire: Donald Trump: 52% Hillary Clinton: 41% #EleccionesEEUU #ElectionDay https://t.co/uhnyqN3ZuC
UniversityWatc1|_HankRearden|0.2732|0.0|0.905|0.095|"RT @_HankRearden: I live in deep blue Boulder, in probably the bluest neighborhood. I've seen literally two Hillary signs total. The energy"
cmpnwtr|FrankLuntz|0.6369|0.0|0.733|0.267|"RT @FrankLuntz: The numbers I'm getting now suggest a nationwide turnout that strongly favors Hillary.And if Hillary does well, so will d"
elllaavalentine|Cj15ive|0.0|0.0|1.0|0.0|RT @Cj15ive: if you vote for Hillary unfollow me
luminouslylit|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: This one's for you, Hillary. https://t.co/KtzpIpSziO"
luminouslylit|twitter|0.0|0.0|1.0|0.0|"RT @HillaryClinton: This one's for you, Hillary. https://t.co/KtzpIpSziO"
jeanne_tall|Caveman2743|0.4466|0.0|0.827|0.173|"RT @Caveman2743: RED ALERT: On Eve of Election, Benghazi BOMBSHELL Rains Down on Hillary https://t.co/rGox20vXgM"
jeanne_tall|conservativetribune|0.4466|0.0|0.827|0.173|"RT @Caveman2743: RED ALERT: On Eve of Election, Benghazi BOMBSHELL Rains Down on Hillary https://t.co/rGox20vXgM"
berkleyparton|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
SLovelace76|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
SLovelace76|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
lewlove123|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
lewlove123|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
emyjeannn|philsadelphia|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
emyjeannn|twitter|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
freerepublican|michelekirkBPR|0.5106|0.0|0.829|0.171|RT @michelekirkBPR: Pro-Hillary rapper marches thousands of fans to Chicago voting booth after free concert https://t.co/j1iz3idvDL https:/
freerepublican|bizpacreview|0.5106|0.0|0.829|0.171|RT @michelekirkBPR: Pro-Hillary rapper marches thousands of fans to Chicago voting booth after free concert https://t.co/j1iz3idvDL https:/
ksootaeho|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
ksootaeho|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
emilyb77|catoletters|-0.5859|0.213|0.787|0.0|RT @catoletters: She has long  history of collaboration with Neocon Warmongers  on foreign policy https://t.co/sSHaBRnVUV
emilyb77|theintercept|-0.5859|0.213|0.787|0.0|RT @catoletters: She has long  history of collaboration with Neocon Warmongers  on foreign policy https://t.co/sSHaBRnVUV
ChiefMya|haylealsina|-0.8934|0.342|0.588|0.07|@haylealsina shit I'd rather Hillary . Because trump just hell naw . He racist af . Like tf ... And if he become president it's over for us
ElisaDonahue|JackPosobiec|-0.2023|0.141|0.859|0.0|RT @JackPosobiec: LIVE on #Periscope: Hillary Workers Intimidate Voters in Philly https://t.co/u9aM89xnPY
ElisaDonahue|periscope|-0.2023|0.141|0.859|0.0|RT @JackPosobiec: LIVE on #Periscope: Hillary Workers Intimidate Voters in Philly https://t.co/u9aM89xnPY
InsaneTrvpper|kiingdarry|0.6249|0.102|0.665|0.232|"RT @kiingdarry: all y'all saying y'all not voting b/c y'all don't believe in Hillary nor Trump, if trump wins Y'ALL BETTER NOT COMPLAIN ABO"
eridani99|donnajherren|-0.6597|0.188|0.812|0.0|"RT @donnajherren: My other kid's speech teacher told her Hillary Clinton has people murdered.Me: Only if they need killing, pumpkin.(YE"
sinncityx|localblactivist|0.0|0.0|1.0|0.0|RT @localblactivist: This correlates to the many instances Trump has pointed out Hillarys war-mongering activities and wall street ties.
kirkbull|dale_bernadette|-0.4574|0.166|0.834|0.0|RT @dale_bernadette: @seanhannity Pennsylvania voters complained of their vote 2 Trump wld switch to Hillary. Frauding again?!
AmBricholas|angryblackhoemo|-0.3595|0.122|0.878|0.0|"RT @angryblackhoemo: white liberals: ""I'm voting for Clinton to stop Trump's racism!""Black people: *lists out ways Hillary's also a racis"
breelieber|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
breelieber|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
dlott1989|hillary_gibble|0.6467|0.0|0.318|0.682|@hillary_gibble @DineshDSouza wonderful!!
tdotsavage00|twitter|0.8225|0.0|0.591|0.409|When u wanted hillary to win but Trump might actually win #distewmuch #andimeanthat https://t.co/TI9ktXGH4N
LDrogosPhD|BitchestheCat|0.0|0.0|1.0|0.0|"RT @BitchestheCat: Every time a state gets called for Hillary, I'm doing a line of catnip. #ElectionDay https://t.co/kuqCiIhtLb"
LDrogosPhD|twitter|0.0|0.0|1.0|0.0|"RT @BitchestheCat: Every time a state gets called for Hillary, I'm doing a line of catnip. #ElectionDay https://t.co/kuqCiIhtLb"
tjcurtis13|AfroGumOfficiaI|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
tjcurtis13|twitter|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
RichardW_1943|DrMartyFox|-0.296|0.121|0.879|0.0|RT @DrMartyFox: #ImVotingBecause We Must Stop DUAL #JUSTICEWhere #Deplorables Must Follow The #RuleOfLawWhile #Hillary &amp; Her Cronies
LayLay_65|MrCouture|0.0|0.0|1.0|0.0|RT @MrCouture: Some of y'all didn't vote but y'all gon be the first ones in line for them Hillary 12's tomorrow!  #ImWithHER https://t.co
LayLay_65|t|0.0|0.0|1.0|0.0|RT @MrCouture: Some of y'all didn't vote but y'all gon be the first ones in line for them Hillary 12's tomorrow!  #ImWithHER https://t.co
CeneJimmy|marwannafuq|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
CeneJimmy|twitter|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
AlishaMichajl|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
pappukepapa|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
amswank|micahwavee|0.802|0.0|0.647|0.353|RT @micahwavee: I think Hillary &amp; Trump supporters alike can at least agree that Branstad needs to go lol.
_JTovar|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
da_realPJay|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
da_realPJay|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
moyankeefan|cascamike|0.0|0.0|1.0|0.0|RT @cascamike: couple of bernie bros voting to put hillary clinton in the white house. https://t.co/2fWUNgWQzK
moyankeefan|twitter|0.0|0.0|1.0|0.0|RT @cascamike: couple of bernie bros voting to put hillary clinton in the white house. https://t.co/2fWUNgWQzK
ayala_joa|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
aeriaIview|hyejenog|0.0|0.0|1.0|0.0|@hyejenog hillary will END him
Ih8heels|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
SulkingWriter|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
SulkingWriter|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
erneststewart6|TruthFeedNews|0.4574|0.16|0.566|0.273|"RT @TruthFeedNews: WOW! HILLARY'S NUMBERS HAVE COLLAPSED IN REUTERS ""TURNOUT"" POLL https://t.co/rAjk98P9kt"
erneststewart6|truthfeed|0.4574|0.16|0.566|0.273|"RT @TruthFeedNews: WOW! HILLARY'S NUMBERS HAVE COLLAPSED IN REUTERS ""TURNOUT"" POLL https://t.co/rAjk98P9kt"
mydogken|MichelleRehorka|-0.69|0.257|0.687|0.056|"@MichelleRehorka @cnnbrk and when Hillary loses, the same gonna happen. Any excuse to tear something up and hurt people!"
awe_rare|ollaollu|0.0|0.0|1.0|0.0|"RT @ollaollu: Hillary: 67,223 votes (29.1%)Trump: 154,176 votes (66.8%)LIVE 6:57:09 PM ET"
babyybry|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
babyybry|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
alecialynn|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
alecialynn|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
_jaycheat|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
a_mamii6|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
kf4bef|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
HansVonSell|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
HansVonSell|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
WmScottBlair|FeliciaBGomez|-0.298|0.149|0.744|0.106|"RT @FeliciaBGomez: Translation: ""We just realized that Hillary's LOSING in NC! Quick! Change the rules! Who cares if it's on the actual ele"
24kcrownn|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
24kcrownn|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
lmjaddict|chasemylovex|0.4404|0.0|0.873|0.127|RT @chasemylovex: Y'all better be throwing away these troll ballots after y'all post these pics for RTs and vote for Hillary.
waughbr|seanhannity|0.0|0.0|1.0|0.0|@seanhannity @realDonaldTrump frank lungs just called the election for Hillary?
grimylittleboy|anuscosgrove|0.0|0.0|1.0|0.0|RT @anuscosgrove: im so high i just typed in google is Hillary or Clinton gonna be president
danhancox|politico|-0.5574|0.153|0.847|0.0|Was trying to explain/recall the nasty tone of the Hillary (+ Bill) 08 primary campaign against Obama and found this https://t.co/HgxylIgdsQ
jesylroche|sadgallexi|-0.5106|0.142|0.858|0.0|"RT @sadgallexi: ""Hillary is a liar, listen to me while I parrot things people have been saying for years to sound smart."" https://t.co/sN2A"
jesylroche|t|-0.5106|0.142|0.858|0.0|"RT @sadgallexi: ""Hillary is a liar, listen to me while I parrot things people have been saying for years to sound smart."" https://t.co/sN2A"
brendanoe60|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
perkoflaura|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
perkoflaura|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
Philly4Really|VanityFair|0.0|0.0|1.0|0.0|RT @VanityFair: Sarah Paulson transforms Hillary Clintons e-mails into award-worthy theater https://t.co/Umx1lB7hsQ https://t.co/GntDhkshBz
Philly4Really|vanityfair|0.0|0.0|1.0|0.0|RT @VanityFair: Sarah Paulson transforms Hillary Clintons e-mails into award-worthy theater https://t.co/Umx1lB7hsQ https://t.co/GntDhkshBz
DUKE_NUKEM_69|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
HIzamoron|Scarlett210|-0.765|0.28|0.72|0.0|"RT @Scarlett210: And #Hillary is a self-serving #elitist who'll continue #globalist policies, destroy ur safety&amp; deprive ur kids of a futur"
Koipan23|JordanRae_24|0.0|0.0|1.0|0.0|RT @JordanRae_24: a lot of people are tryna vote for trump but the computers are changin it to Hillary 
SaraVespucci|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
SaraVespucci|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
lookitslyndseyy|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
IAmTayNelson|___DestinyJadai|-0.6739|0.476|0.524|0.0|"RT @___DestinyJadai: ""VOTE HILLARY BITCH""  https://t.co/xVltWc6dU7"
IAmTayNelson|twitter|-0.6739|0.476|0.524|0.0|"RT @___DestinyJadai: ""VOTE HILLARY BITCH""  https://t.co/xVltWc6dU7"
creminsmom|JOHNSONSFOOL|-0.4003|0.119|0.881|0.0|@JOHNSONSFOOL If Hillary worked for a bank (any US Company) &amp;  released Confidential Info.... She is fired.... Fire Hillary .... Vote Trump!
serena_223|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
serena_223|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
_Zakkery_|FreeMemesKids|-0.1695|0.196|0.804|0.0|"RT @FreeMemesKids: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
stumpyyyyyyy|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
crose84|Lisa_JDC|0.0|0.0|1.0|0.0|"RT @Lisa_JDC: If you were in line before the polls close, you have the right to vote. #StayInLine and vote for #hillary #ElectionDay https:"
jamesedgriffin|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
jamesedgriffin|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
LaurynKhleo|mefeater|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
LaurynKhleo|twitter|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
_IHateIgnorance|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
ntamylee|FIirtationship|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
ntamylee|twitter|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
rdonoghue|Spacekatgal|0.5106|0.0|0.875|0.125|"RT @Spacekatgal: CSPAN is passing out free copies of the constitution at Hillary HQ, which is the most C-SPAN thing to do ever. #ImWithHer"
sorrowen|TwitchyTeam|0.296|0.0|0.879|0.121|"RT @TwitchyTeam: Guy Benson shares Hillarys internals via a Dem source, take with grains of salt #ElectionNight https://t.co/BvrwdS5WIh"
sorrowen|twitchy|0.296|0.0|0.879|0.121|"RT @TwitchyTeam: Guy Benson shares Hillarys internals via a Dem source, take with grains of salt #ElectionNight https://t.co/BvrwdS5WIh"
hannah_leeann16|StevannaA|0.3832|0.101|0.71|0.189|RT @StevannaA: It blows my mind that so many Americans who were raised to value honesty are completely ignoring the fact that Hillary CANNO
JJManring|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
JJManring|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
Rich_893|billmaher|-0.8753|0.382|0.574|0.044|"RT @billmaher: Pls vote for Hillary today. Even if you don't like her, its necessary to block a dangerous lunatic ultimate power. #ThisTime"
POLITICAL_Jeff|mitchellvii|-0.7645|0.32|0.68|0.0|"RT @mitchellvii: Based upon exits, voters very unhappy with big money corruption.  That's bad for Hillary."
EmehDR|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
EmehDR|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
samkrenz_|billmaher|-0.8753|0.382|0.574|0.044|"RT @billmaher: Pls vote for Hillary today. Even if you don't like her, its necessary to block a dangerous lunatic ultimate power. #ThisTime"
_tierrrraaaa|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_tierrrraaaa|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Khaleesi_Hodan|TheDailyShow|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
Khaleesi_Hodan|cc|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
demar19511|linkis|0.5719|0.0|0.764|0.236|Pat Buchanan Says The Country Will &amp;#8216;Not Be United&amp;#8217; If Hillary Wins: https://t.co/WtIwOcQxrM
d6sty|PzFee|0.4404|0.0|0.873|0.127|RT @PzFee: BREAKING NEWS -- Spongebob shot at Trump rally. He was supporting Hillary Clinton and got shot by Plankton. https://t.co/mU8MRF2
d6sty|t|0.4404|0.0|0.873|0.127|RT @PzFee: BREAKING NEWS -- Spongebob shot at Trump rally. He was supporting Hillary Clinton and got shot by Plankton. https://t.co/mU8MRF2
lilwha13|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
lilwha13|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
the_Jordanrules|Dolo_kd|0.0|0.111|0.777|0.111|RT @Dolo_kd: I'm voting for Hillary Clinton only because she's a strong woman who stood by her husband side after he cheated .. she has cha
carefreegrldom|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
carefreegrldom|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
_DonnyT|giveyouIife|-0.128|0.2|0.8|0.0|RT @giveyouIife: cutting up for Hillary https://t.co/jPUGgWhB8K
_DonnyT|twitter|-0.128|0.2|0.8|0.0|RT @giveyouIife: cutting up for Hillary https://t.co/jPUGgWhB8K
Hardline_Stance|He_Has_Failed|-0.6486|0.306|0.694|0.0|"RT @He_Has_Failed: Hillary Ally Warned She, Dems Could Be Destroyed By Corruption https://t.co/ZO7FCMi8kO https://t.co/X3Gvtjyi16"
Hardline_Stance|dailycaller|-0.6486|0.306|0.694|0.0|"RT @He_Has_Failed: Hillary Ally Warned She, Dems Could Be Destroyed By Corruption https://t.co/ZO7FCMi8kO https://t.co/X3Gvtjyi16"
pacmann007|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
pacmann007|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
lopezzjenn|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
DunkirkDavid|jakerock88|0.7003|0.0|0.746|0.254|@jakerock88 good evening Jake thanks for the follow we need Donald Trump as our president never Hillary @TeamTrump #Election2016
StephanieMitz|FemMajority|0.0|0.0|1.0|0.0|"RT @FemMajority: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https"
TuNaLdO|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
TuNaLdO|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
becky_page_|Kay_wizz1|-0.1182|0.1|0.819|0.082|"RT @Kay_wizz1: But Hillary can't be trusted w her own email account. Which is to me, a lot more important that twitter. Don't @ me https://"
becky_page_||-0.1182|0.1|0.819|0.082|"RT @Kay_wizz1: But Hillary can't be trusted w her own email account. Which is to me, a lot more important that twitter. Don't @ me https://"
kmichelleregus|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
kmichelleregus|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
KeilaCee|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
azdespot|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
azdespot|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
JIndeliclae|brainpicker|-0.6597|0.24|0.702|0.058|"RT @brainpicker: ""Im horrified to watch the bizarre pageant of my nation pretending these two contenders are equivalent."" THIS https://t.c"
JIndeliclae||-0.6597|0.24|0.702|0.058|"RT @brainpicker: ""Im horrified to watch the bizarre pageant of my nation pretending these two contenders are equivalent."" THIS https://t.c"
V_Krassilnikov|foreignpolicy|0.0|0.0|1.0|0.0|The Hillary Clinton Doctrine https://t.co/T3P0Lb7rE3
caleb_330|Avstvn|-0.1695|0.196|0.804|0.0|"RT @Avstvn: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
miraculashton|HillaryClinton|0.6486|0.0|0.819|0.181|"RT @HillaryClinton: ""I believe with all my heart that our best days are still ahead of us, if we reach for them together. Hillary in Phil"
vlenxx|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
vlenxx|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
hotteronline|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
princessmyaxa|Katie__Huang|0.8894|0.0|0.666|0.334|RT @Katie__Huang: FRIENDLY REMINDER THAT IF HILLARY WINS BERNIE WILL BE HEAD OF SENATE BUDGET COMMITTEE IF DEM GET THE MAJORITY!!!!!!
schmerielle|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
schmerielle|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
BryanCusick|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
BryanCusick|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
greggypoo65|xmssweetnessx|0.34|0.192|0.5|0.308|"RT @xmssweetnessx: If Hillary Wins, America Loses  #WTFAmericaIn5Words"
cheyennenicoleg|a_adams23|0.0|0.0|1.0|0.0|RT @a_adams23: How to vote for Hillary Clinton https://t.co/w4pOBMTGPn
cheyennenicoleg|twitter|0.0|0.0|1.0|0.0|RT @a_adams23: How to vote for Hillary Clinton https://t.co/w4pOBMTGPn
TheMinerK|TheFunnyVine|-0.0191|0.097|0.903|0.0|RT @TheFunnyVine: Trump and Hillary will never reach this level  https://t.co/9jl1rDKqj7
TheMinerK|vine|-0.0191|0.097|0.903|0.0|RT @TheFunnyVine: Trump and Hillary will never reach this level  https://t.co/9jl1rDKqj7
emileemaeeeh|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
marianperales_|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
marianperales_|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Ammirzi|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Ammirzi|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
willOBell|AmiriKing|0.0|0.0|1.0|0.0|RT @AmiriKing: Idea:Split the U.S. in half.Dems get one side.Reps get one side.Hillary runs your lives.Trump leads ours.#Clinto
ryncarnate|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
CharliseAnne|ClarenceJWhite|0.0|0.069|0.863|0.069|RT @ClarenceJWhite: I feel like Trump &amp; Hillary are two divorced parents fighting over custody of us but we kinda just wanna go live with g
jamieefoster|DanaSchwartzzz|0.6249|0.075|0.712|0.214|RT @DanaSchwartzzz: Dear lord if Hillary Clinton wins I'll read a book before bed and stop tweeting so much and give more to the homeless a
Nikki_Bitchhh|ShineVista|0.3616|0.148|0.608|0.243|"RT @ShineVista: Prediction: Hillary Clinton wins election, Donald Trump doesn't concede. America riots, &amp; people die. Market crashes. Haram"
VeriteGrace|youtube|0.0|0.0|1.0|0.0|Julian Assange Drops BOMBSHELL on Hillary Clinton https://t.co/lUQVzgEmhQ
enamoramiento1|lizcgoodwin|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
enamoramiento1|twitter|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
erythingistaken|cykelly1718|0.6808|0.0|0.741|0.259|"@cykelly1718 @hindman_ben @HillaryClinton I am in Diamond Business,I just happened to care for poor,I am a millionair.I still think HILLARY."
JerryGrinstead|ed_hooley|-0.8769|0.404|0.485|0.111|RT @ed_hooley: HILLARY'S VP TIM KAINE REFUSED TO HELP ME. DAUGHTER KILLED BY ILLEGAL IMMIGRANT #ElectionDay #ElectionNight #RAW https://t.
JerryGrinstead||-0.8769|0.404|0.485|0.111|RT @ed_hooley: HILLARY'S VP TIM KAINE REFUSED TO HELP ME. DAUGHTER KILLED BY ILLEGAL IMMIGRANT #ElectionDay #ElectionNight #RAW https://t.
pplenkie|JackPosobiec|-0.8668|0.52|0.48|0.0|RT @JackPosobiec: SHOCK VIDEO: Hillary Workers Violently Threaten Voters in W Philly https://t.co/J76EcwbZhZ
pplenkie|periscope|-0.8668|0.52|0.48|0.0|RT @JackPosobiec: SHOCK VIDEO: Hillary Workers Violently Threaten Voters in W Philly https://t.co/J76EcwbZhZ
edenrathore|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
edenrathore|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
brandoniii12|piratejeffrey|-0.5562|0.253|0.625|0.121|RT @piratejeffrey: Whoa this kinda blows your mind! Brutally honest story of the feminist Hillary Rodham we desperately need...  https:/
brandoniii12||-0.5562|0.253|0.625|0.121|RT @piratejeffrey: Whoa this kinda blows your mind! Brutally honest story of the feminist Hillary Rodham we desperately need...  https:/
JulieCTaylor|worldnetdaily|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
JulieCTaylor|wnd|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
SuzieQt154320|Pamela_Moore13|-0.5386|0.267|0.595|0.138|RT @Pamela_Moore13: Man PROVES software stole votes in ALL 'Hillary won' counties! DNC rigged elections!Voter Fraud is Real! https://t.co
SuzieQt154320|t|-0.5386|0.267|0.595|0.138|RT @Pamela_Moore13: Man PROVES software stole votes in ALL 'Hillary won' counties! DNC rigged elections!Voter Fraud is Real! https://t.co
stabley2|MadelnCanada|0.0|0.0|1.0|0.0|@MadelnCanada Hillary*
alpha_joe86|Things4Guys|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
alpha_joe86|twitter|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
cesarleeon1|Pasion_Basket|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
cesarleeon1|twitter|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
sergiocancelo|Pasion_Basket|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
sergiocancelo|twitter|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
everydaydolans|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
babybookay|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
babybookay|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Rayaa001|PoppinAssMia|-0.4023|0.311|0.689|0.0|RT @PoppinAssMia: I don't trust Hillary or Trump 
JJCobb1_|Raven_Babby_|0.0|0.0|1.0|0.0|"RT @Raven_Babby_: I'm behind Obama, &amp; he's behind Hillary "
brizeemode|DarriusKV|0.0772|0.0|0.885|0.115|"RT @DarriusKV: Vote for who you want, vote for Hillary https://t.co/oxGyhowtEt"
brizeemode|twitter|0.0772|0.0|0.885|0.115|"RT @DarriusKV: Vote for who you want, vote for Hillary https://t.co/oxGyhowtEt"
Santy0722|TrashvisScott|0.5719|0.0|0.764|0.236|RT @TrashvisScott: if Hillary wins I'll PayPal $1 to everyone who RTs this 
heeidi___|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
heeidi___|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
gerry_dankowski|PrisonPlanet|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
gerry_dankowski|pittsburgh|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
annamurack22|CloydRivers|0.0|0.0|1.0|0.0|RT @CloydRivers: Im not against a woman bein President. Im just against that woman bein Hillary Clinton. Merica.
pithypisces|jb19tele|0.0|0.0|1.0|0.0|RT @jb19tele: James O'Keefe Files FEC Suit Against Hillary Clinton - Breitbart https://t.co/7QH8MugNYM via @BreitbartNews
pithypisces|linkis|0.0|0.0|1.0|0.0|RT @jb19tele: James O'Keefe Files FEC Suit Against Hillary Clinton - Breitbart https://t.co/7QH8MugNYM via @BreitbartNews
_s0ire|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_s0ire|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
KuldeepRaina15|BDUTT|0.4019|0.0|0.886|0.114|RT @BDUTT: Live from the Glass Ceiling I bet Hillary Clinton Will Smash tonight. The venue of her Victory Party. Facebook Live https://t.co
KuldeepRaina15|t|0.4019|0.0|0.886|0.114|RT @BDUTT: Live from the Glass Ceiling I bet Hillary Clinton Will Smash tonight. The venue of her Victory Party. Facebook Live https://t.co
mennahamed8|TheAdly|-0.1027|0.065|0.935|0.0|"RT @TheAdly: #Hillary or #Trump, America will make history today. Either the first female president, or the first mentally challenged one."
brockjamiedave|LeighPatrick|0.0|0.0|1.0|0.0|"RT @LeighPatrick: Given the reports flooding in nationwide, you either vote Hillary or the machine votes Hillary for you. #Corruption #elec"
ChuckNellis|SneakyBlackDog|0.0|0.0|1.0|0.0|@SneakyBlackDog So he's conceding Hillary wins...
Labeez_|twitter|-0.3182|0.195|0.7|0.105|"Me when Hillary ignored the cries for help from Ambassador Stevens, Sean Smith, Glen Doherty, &amp; Tyrone Woods, &amp; let https://t.co/2kcIvSNsUw"
leancar2010|johnauthers|0.5256|0.0|0.861|0.139|RT @johnauthers: Forex markets now betting more confidently on Hillary. Dollar continuing to fall vs Mexican peso. Brexit II or right secon
ShrekLover6969|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
DaveyHo69|_nswerhunmain_|-0.5216|0.195|0.805|0.0|RT @_nswerhunmain_: Hillary can't protect FOUR Americans in Benghazi... How is she going to protect the whole country? #TrumpPence16  #Ele
BradTurner39|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
Kayx2__|chasemylovex|-0.3586|0.127|0.873|0.0|"RT @chasemylovex: no, Hillary is not the ""ideal candidate"" but we still gonna vote for her tho... and we'll deal with sis later, ya hear me"
Sensei_Ensell|KayzoMusic|0.765|0.0|0.68|0.32|RT @KayzoMusic: If Hillary Clinton wins I hope she comes out for her victory speech to jotaro.
BeachAddict80|FoxBusiness|0.5859|0.0|0.863|0.137|"RT @FoxBusiness: .@ktmcfarland: ""If [#Hillary] does win, she is not going to be able to govern. She has so much baggage, she is so corrupt."
RuiMalbreezyDBz|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Ayoobray_|GIRLHEFUNNY|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
Ayoobray_|twitter|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
Adriana_Lopez87|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
Adriana_Lopez87|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
OneTrump4All|ppetrov5|0.0|0.0|1.0|0.0|"RT @ppetrov5: Hillary Clinton and her campaign met with prioritiesUSA, which is against the law. #PodestaEmails35 #wikileaks #fbi https://t"
OneTrump4All||0.0|0.0|1.0|0.0|"RT @ppetrov5: Hillary Clinton and her campaign met with prioritiesUSA, which is against the law. #PodestaEmails35 #wikileaks #fbi https://t"
reignonu|kt_taylor17|0.3612|0.0|0.898|0.102|"RT @kt_taylor17: when i wake up in the morning, im praying thata) hillary will be president b) there'll be a steaming plate of katsu next"
babycilla_|RiRiHumor|0.0|0.0|1.0|0.0|RT @RiRiHumor: Rihanna wearing a shirt of a picture of herself wearing a Hillary Clinton shirt. She's with HER! #ElectionDay https://t.co/X
babycilla_|linkedin|0.0|0.0|1.0|0.0|RT @RiRiHumor: Rihanna wearing a shirt of a picture of herself wearing a Hillary Clinton shirt. She's with HER! #ElectionDay https://t.co/X
gaabiwalsh|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
DeeDub8|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
blueefoxxx|Ekatherene|0.0|0.0|1.0|0.0|"RT @Ekatherene: @mitchellvii @MarianneHaran Las Vegas has Hillary down by 7% , last night she was down 5%...."
JazmineMejia14|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
JazmineMejia14|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
kirstenstauffe1|LondraPolitics|0.0|0.0|1.0|0.0|"RT @LondraPolitics: According to the Turkish media funded by Erdogan, here is the first #ElectionNight exit poll results;Hillary: 20%Tru"
jsrroger|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @Slate @votecastr @LilSteelerGirl @DebAlwaystrump @Kerri1111 TRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLID
rayven_alexa|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
rayven_alexa|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
CCrusherP|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
supbrea|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
JakaylaLovesYou|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
JakaylaLovesYou|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
__damnitsdiaaa|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
__damnitsdiaaa|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
BackmanMegan|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
BackmanMegan|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
HerbApproach|theweedblog|0.0|0.0|1.0|0.0|Why Hillary Clinton Could be More Than the First https://t.co/22pBl7AV3J #Ending_Marijuana_Prohibition #election_2016 #hillary_clinton
Jackiie_Salinas|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
LUSTlG|open|-0.6956|0.345|0.655|0.0|#NowPlaying FDT but also fuck hillary too by YG  https://t.co/g4DgIPWVyV
gracieeisabelle|haquimo_|0.5719|0.0|0.619|0.381|RT @haquimo_: Me if Hillary wins https://t.co/RPPuzbJddB
gracieeisabelle|twitter|0.5719|0.0|0.619|0.381|RT @haquimo_: Me if Hillary wins https://t.co/RPPuzbJddB
gutierrezy14|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
gutierrezy14|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Erictrevisan1|RobinDavani|-0.8941|0.339|0.661|0.0|RT @RobinDavani: @celestemc @CNNPolitics MORE VOTER FRAUD IN DURHAM COUNTY NC! 90 MINUTE EXTENSION TO CAST FRAUDULENT VOTES FOR HILLARY ALL
Rayy1567|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
ShuB0x|Eliza24___|0.5719|0.0|0.837|0.163|"RT @Eliza24___: Hillary won Kentucky. We are still waiting on the results from Mcdonald's, Wendy's, Burger King and Taco Bell."
Jarret_Stanton|WesVengeance7|0.296|0.0|0.891|0.109|RT @WesVengeance7: The joke is on Hillary if she wins.She'll have to sit at the desk Monica sat under.
crescentegus|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
crescentegus|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
scuttigirl|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
scuttigirl|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
bridgetmarian|ImDaddysAngel|-0.5106|0.121|0.879|0.0|RT @ImDaddysAngel: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote f
MarcoAD80|thedoubleb|0.1027|0.242|0.549|0.209|"@thedoubleb wow, dirty tricks. Hickey is a Republican who opposes Hillary. Vote Democrat @MaraWElliott"
DiSwanson77|andersonDrLJA|-0.8122|0.286|0.714|0.0|RT @andersonDrLJA: #Crooked HILLARY HERSELF HAS SAID No One Is To Big to be Prosecuted &amp; Sent to Prison SO BE IT! #HillaryForPrison2016 htt
_NoFilter_|_ShowNoLovee|0.0|0.0|1.0|0.0|@_ShowNoLovee trump and Hillary 
VeeLo_Greene|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
gibsonnbecca|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
gibsonnbecca|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
jonnothorsley|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
jonnothorsley|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
rowanevejones|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
lvcymiller|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
lvcymiller|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
IM_extrAVAgant|Inc|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
IM_extrAVAgant|t|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
bearoserod|BuzzFeedNews|-0.7028|0.271|0.729|0.0|"RT @BuzzFeedNews: 29 Most WTF Moments Of The Election: Hillary's Trump ""Joke"" #ElectionDay https://t.co/PNF7xkBxgB"
bearoserod|twitter|-0.7028|0.271|0.729|0.0|"RT @BuzzFeedNews: 29 Most WTF Moments Of The Election: Hillary's Trump ""Joke"" #ElectionDay https://t.co/PNF7xkBxgB"
Winky2124|_cam_white_|0.128|0.088|0.805|0.107|"RT @_cam_white_: When Hillary was asked about the American lives lost in Benghazi her response was ""What does it matter"". Vote Wisely #TRUM"
gocoo|TheVampsJames|0.0|0.0|1.0|0.0|"RT @TheVampsJames: 2 years ago in radio 2, Tris and I were walking out and we saw Hillary Clinton. She said to us 'you're the vamps right?'"
adorehails|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
adorehails|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
Katiecook55|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
Katiecook55|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
helovedmemore|dyanjae|0.1012|0.104|0.776|0.121|RT @dyanjae: @mitchellvii Doug Schoen said internal FL Hispanic vote is around 50-30+ &amp; if true not good for Hillary.
Skydawgy1|TomiLahren|0.4717|0.0|0.861|0.139|RT @TomiLahren: If you're not voting for Trump don't you dare bitch when we get Hillary. Real talk. #MAGA #ElectionDay
GuapoDaGawd|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
GuapoDaGawd|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Joan_Ripolles|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  (cont) https://t.co/y61yMeEMLE
Joan_Ripolles|twitlonger|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  (cont) https://t.co/y61yMeEMLE
rawcurrent|bendandSNAPPER|0.0|0.0|1.0|0.0|RT @bendandSNAPPER: Find someone who looks at you the way Hillary looks at balloons. https://t.co/Lmyu5HDvjk
rawcurrent|twitter|0.0|0.0|1.0|0.0|RT @bendandSNAPPER: Find someone who looks at you the way Hillary looks at balloons. https://t.co/Lmyu5HDvjk
miraculashton|HillaryClinton|0.1421|0.12|0.783|0.098|"RT @HillaryClinton: ""We dont want to shrink the vision of this country. We want to keep expanding it. Hillary"
171312Joe|kevvgallagher|0.7717|0.1|0.592|0.308|"RT @kevvgallagher: Lmao if you're a Republican and get mad when Hillary wins, maybe you should've supported one of the other 16 options. It"
CloverOG|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
CloverOG|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
HammLogan|twitter|-0.3612|0.161|0.839|0.0|you know Hillary was fighting off having a seizure while trying to stay still https://t.co/ZRztImwiAs
bringitbri_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
GagAlexFrance|musicnews_facts|0.4404|0.0|0.873|0.127|"RT @musicnews_facts: Trump supporters are calling out Hillary Clinton and Lady Gaga for wearing this ""Nazi Hitler"" uniform... When it's Mic"
DanTillotson|HaroldItz|0.4926|0.0|0.856|0.144|@HaroldItz He we go then Harold. Let's hope that filthy sleaze bag gets a spanking. Go Hillary! Is the scotch out?
kingnessaa|JOHNSONSFOOL|0.7579|0.0|0.727|0.273|"RT @JOHNSONSFOOL: you still have time, please please go vote for hillary, she's the better option for you &amp; the youths future #ElectionNigh"
BusinessNews40|marketwatch|0.0|0.0|1.0|0.0|Unlikely fashion icon Hillary Clinton is bringing back the pantsuit https://t.co/gycJZFnXTq #Business https://t.co/SzeLp351MU
SandraKennett1|LouDobbs|-0.7574|0.372|0.544|0.083|"@LouDobbs Hillary isn't well liked by people, while Donald Trump is loved by people, but not well liked by the biased MSM."
MeganNemec|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
MeganNemec|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
colewells1001|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
SomeGuysCat|JohnFromCranber|0.6739|0.0|0.835|0.165|RT @JohnFromCranber: It's All About Turnout. Typically Only About 1/2 Vote. If All the Folks who Prefer Trump Over Hillary Vote - WE WIN IN
Stairmaster_|SluttySam2|-0.7003|0.286|0.611|0.103|"RT @SluttySam2: ""I hate hillary""""That means you support sexual assault and racism""""...No, that's not what that means at all"""
Max2Min|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Max2Min|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
haddynuff|StopStopHillary|0.0|0.0|1.0|0.0|RT @StopStopHillary: FIRST POLLS FOR KENTUCKY TRUMP 78%HILLARY 18%
buteraftommo|musicnews_facts|0.0|0.0|1.0|0.0|RT @musicnews_facts: Lady Gaga spoke at a Hillary Clinton rally tonight wearing a Michael Jackson military attire. https://t.co/rYJUL805Ae
buteraftommo|twitter|0.0|0.0|1.0|0.0|RT @musicnews_facts: Lady Gaga spoke at a Hillary Clinton rally tonight wearing a Michael Jackson military attire. https://t.co/rYJUL805Ae
_life_as_tay|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
_life_as_tay|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
aislam_|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
JoeRiggs10|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
max_weidman|WesVengeance7|0.296|0.0|0.891|0.109|RT @WesVengeance7: The joke is on Hillary if she wins.She'll have to sit at the desk Monica sat under.
JustGoForIt|skyhookmike|-0.7254|0.272|0.728|0.0|RT @skyhookmike:  Because no REAL man WANTED that FILTHY MOUTH on their DI#%! Madonna Won't Honor Promise to Fellate Hillary Voter https:/
JustGoForIt||-0.7254|0.272|0.728|0.0|RT @skyhookmike:  Because no REAL man WANTED that FILTHY MOUTH on their DI#%! Madonna Won't Honor Promise to Fellate Hillary Voter https:/
helghast_chen|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
helghast_chen|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
sameoldsxlena|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
sameoldsxlena|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
ftdbev|DavidCornDC|0.0|0.0|1.0|0.0|RT @DavidCornDC: Where Hillary Clinton will declare victory or....something else. https://t.co/4b82Lt4UGB
ftdbev|twitter|0.0|0.0|1.0|0.0|RT @DavidCornDC: Where Hillary Clinton will declare victory or....something else. https://t.co/4b82Lt4UGB
Krakenpodcast|twitter|0.3291|0.0|0.885|0.115|googoo gaga. ken loves barbie BUT barbie is hillary. my takes would justify george r r martin's premature demise an https://t.co/sqFobr8wQr
nwjerseyliz|CNN|0.4019|0.0|0.863|0.137|RT @CNN: Women across the nation are wearing pantsuits on #ElectionDay in support of Hillary Clinton https://t.co/TN3TeGDuDi #Pantsuitnatio
nwjerseyliz|cnn|0.4019|0.0|0.863|0.137|RT @CNN: Women across the nation are wearing pantsuits on #ElectionDay in support of Hillary Clinton https://t.co/TN3TeGDuDi #Pantsuitnatio
JeonsRoyalty|SuelovesBts|-0.1027|0.123|0.877|0.0|@SuelovesBts @Iovespell They even got a Hillary one idk what's going on
kittycatbaty|DonaldJTrumpJr|0.5719|0.0|0.73|0.27|"RT @DonaldJTrumpJr: Sean Hannity: If Hillary wins, you own it https://t.co/Wo8k89T7s9"
kittycatbaty|video|0.5719|0.0|0.73|0.27|"RT @DonaldJTrumpJr: Sean Hannity: If Hillary wins, you own it https://t.co/Wo8k89T7s9"
murgaloo|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
_Byethai|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_Byethai|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
bistrogal2|twitter|0.5599|0.0|0.859|0.141|"PLEASE EVERYONE.GET OUT &amp; VOTE FOR TRUMP! EVEN IF YOU HAVE A COLD, APPT - ANY REASON, JUST GET OUT &amp; VOTE! DRAIN TH https://t.co/Z7UKiWzkHL"
shxmvllnv|vibeeeez|-0.5574|0.261|0.739|0.0|RT @vibeeeez: prediction: Hillary Clinton is our next present &amp; everyone is shocked Trump lost
Freedom61815022|gs777gs777|-0.893|0.4|0.6|0.0|RT @gs777gs777: I have not seen ONE REPORT of voter fraud by Republicans ! Disgusting dirty campaign by Hillary Clinton ! https://t.co/Q7B0
Freedom61815022|t|-0.893|0.4|0.6|0.0|RT @gs777gs777: I have not seen ONE REPORT of voter fraud by Republicans ! Disgusting dirty campaign by Hillary Clinton ! https://t.co/Q7B0
FirstNameMiaa|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
FirstNameMiaa|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
270Strategies|MarlonDMarshall|0.0|0.0|1.0|0.0|Check out 270's @MarlonDMarshall and @mansara in Hillary's #MannequinChallenge! https://t.co/OQPhnADGlG
270Strategies|twitter|0.0|0.0|1.0|0.0|Check out 270's @MarlonDMarshall and @mansara in Hillary's #MannequinChallenge! https://t.co/OQPhnADGlG
j_taylor_b|brittanymacik|0.7506|0.0|0.652|0.348|RT @brittanymacik: All in favor of Texas seceding from the US if Hillary wins
FrannieC_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
focused_4|Chico_Mills|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
focused_4|twitter|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
clintonchineduc|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana 0.6% reporting TRUMP 69.8% | Hillary 26.4%  massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Elect
macamaw61|chasin_dwight|0.4019|0.088|0.749|0.163|RT @chasin_dwight: #TheFive If Hillary wins I can cancel cable. Will not be able to turn TV on for 4 years
beltranaminta|HaskelBiz|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
beltranaminta|twitter|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
girlnamedjon|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
revsaint08|drewwyatt|-0.5216|0.151|0.849|0.0|RT @drewwyatt: Hillary Campaign Paid Rioters 2 Burn The American Flag @ Trump Rally.You Can't Love Our Country &amp; Justify Voting 4 Her.
jaybabyy_89|chasemylovex|-0.3586|0.127|0.873|0.0|"RT @chasemylovex: no, Hillary is not the ""ideal candidate"" but we still gonna vote for her tho... and we'll deal with sis later, ya hear me"
goodkidgouth|azitatoprahman|0.0|0.0|1.0|0.0|@azitatoprahman did you just assume Hillary's gender
MollyQuilitzsch|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
MollyQuilitzsch|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
EileenPereira_|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
EileenPereira_|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
BrookeSeagrave|FIirtationship|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
BrookeSeagrave|twitter|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
JasonDunn67|PizzaPartyBen|0.0|0.0|1.0|0.0|"RT @PizzaPartyBen: Hillary Clinton's mentor was a leader in the KKK, actually #MyVote2016 #ElectionDay #Voted #TuesdayMotivation https://"
JasonDunn67||0.0|0.0|1.0|0.0|"RT @PizzaPartyBen: Hillary Clinton's mentor was a leader in the KKK, actually #MyVote2016 #ElectionDay #Voted #TuesdayMotivation https://"
frogopera|twitter|0.0258|0.107|0.782|0.111|"""thousands of people are flocking to susan b. anthony's grave in memory of her movement and in support of hillary"" https://t.co/n6Q1B7NZc4"
therealmofnay|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
therealmofnay|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Magical_Grrl|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
Magical_Grrl|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
ohmyswift1213|vibeeeez|-0.5574|0.261|0.739|0.0|RT @vibeeeez: prediction: Hillary Clinton is our next present &amp; everyone is shocked Trump lost
mllnola|DrThomasPaul|0.6114|0.0|0.81|0.19|RT @DrThomasPaul: Happy about this #LGBT/#LGBTQ for anyone who thinks #Hillary is for #gays? Think again!She's financing #murders.#gayhttp
Ssmfarley777|Abutbul9|-0.4767|0.194|0.806|0.0|RT @Abutbul9: Breaking: Hillary Clintons $20 Million Obama Bribe To Become US Secretary Of State Leaked By FBI https://t.co/MIJecsJEP3
Ssmfarley777|endingthefed|-0.4767|0.194|0.806|0.0|RT @Abutbul9: Breaking: Hillary Clintons $20 Million Obama Bribe To Become US Secretary Of State Leaked By FBI https://t.co/MIJecsJEP3
tamaraleighllc|JoeyArnoldVN|0.0|0.0|1.0|0.0|RT @JoeyArnoldVN: GO VOTE TODAY TRUMP HILLARY CLINTON#ExitPoll#iVoted#myVote2016#ElectionDay#VoteJSA#Poll#WTFAmericaIn5Words#DolanT
mr_inkcognito|DontTread_2nd|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
mr_inkcognito|twitter|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
KC__xballoutx|VinePhilly|0.0772|0.0|0.794|0.206|RT @VinePhilly: Hillary Mannequin Challenge https://t.co/NqRLzIcUqN
KC__xballoutx|twitter|0.0772|0.0|0.794|0.206|RT @VinePhilly: Hillary Mannequin Challenge https://t.co/NqRLzIcUqN
Tehpanga|slayinglooks|0.0|0.0|1.0|0.0|RT @slayinglooks: Will Hillary make pants suits mandatory?Will Trump build a wall on Mexicos border?   Find out tomorrow on the season
Graysun182|ianbrink24|-0.7269|0.337|0.663|0.0|RT @ianbrink24: Hillary Clinton's the type of person to hide the cure for cancer.
katgal2|BritsForHill|0.2323|0.101|0.759|0.14|RT @BritsForHill: PLEASE don't assume #Hillary victory is guaranteed...we made that mistake with Brexit. Go out and TAKE IT! #nevertrump
dejean76|gerfingerpoken|0.0|0.0|1.0|0.0|"RT @gerfingerpoken: Trump Defends Life, Hillary Defends #PartialBirthAbortion - Flopping Aces - https://t.co/boHSpqQIqN #MAGA https://t.co/"
dejean76|floppingaces|0.0|0.0|1.0|0.0|"RT @gerfingerpoken: Trump Defends Life, Hillary Defends #PartialBirthAbortion - Flopping Aces - https://t.co/boHSpqQIqN #MAGA https://t.co/"
Tropicblasiann|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Tropicblasiann|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
peaceoutanddab|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
imbeccajett|xD1v1ne|-0.0772|0.337|0.361|0.301|@xD1v1ne @tha_macey Lies. Like Hillary.
SupaKawaiiLexi|ScienceTrash|0.4201|0.0|0.877|0.123|"@ScienceTrash But it still has to go through Congress. I'm not for Trump, or Hillary. So I agree with what you're saying."
VilleSZN|JayeNick_|-0.5719|0.236|0.764|0.0|RT @JayeNick_: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/dpWCWHwHhw
VilleSZN|twitter|-0.5719|0.236|0.764|0.0|RT @JayeNick_: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/dpWCWHwHhw
rtoberl|barb2939|-0.296|0.095|0.905|0.0|RT @barb2939: @magnifier661 @johnpodesta No wonder Hillary moved billion of her money to bank in Quter a few Saturday mornings ago. Or was
blkshirtfan|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
iIoveharry|yvezayntIaurent|-0.5423|0.22|0.78|0.0|"RT @yvezayntIaurent: white person: idk whos worse: hillary or trumplgbtq, women, black people, immigrants, muslims: trump iswhite pers"
M3l3ah|tbscott2|0.5719|0.0|0.684|0.316|RT @tbscott2: If Hillary wins I'm moving to Canada 
bryceMartian54|memetribute|-0.1695|0.186|0.814|0.0|"RT @memetribute: We don't want Trump, we don't want Hillary, we just want Cory back in the house #ElectionDay"
kayy_ash|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
mikedanzar|Jess_P_7385|0.68|0.0|0.728|0.272|RT @Jess_P_7385: If anyone thinks about voting for #Hillary please consider this cute little ducks opinion!#TrumpPence16 #MakeAmericaGreatA
Make_Me_Smil3|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Make_Me_Smil3|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
StevenRuizok|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
StevenRuizok|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
ArthurRFagundes|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
ArthurRFagundes|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
trnichols12|t_howay02|0.6486|0.0|0.675|0.325|RT @t_howay02: Hillary's trash I just don't get why you all like her lol
SmitaRanjit|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
SmitaRanjit|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
JanDupuy|GovMikeHuckabee|0.0|0.0|1.0|0.0|"RT @GovMikeHuckabee: State Dept says it takes 5 yrs to review 31,000 Hillary emails. Let Comey do it!  He can review 650,000 in 1 week!  ht"
vaaaaalarie|DaiIyRap|0.0772|0.0|0.86|0.14|RT @DaiIyRap: Hillary Clinton doing the Mannequin Challenge https://t.co/yZXFZ1hNrn
vaaaaalarie|twitter|0.0772|0.0|0.86|0.14|RT @DaiIyRap: Hillary Clinton doing the Mannequin Challenge https://t.co/yZXFZ1hNrn
lovehope|theGrio|0.4019|0.0|0.87|0.13|RT @theGrio: #Beyonc made one last ditch effort for voters to support #HillaryClinton in this Tidal PSA: https://t.co/GSJe9BqP12 https://t
lovehope|thegrio|0.4019|0.0|0.87|0.13|RT @theGrio: #Beyonc made one last ditch effort for voters to support #HillaryClinton in this Tidal PSA: https://t.co/GSJe9BqP12 https://t
octavenduh|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
octavenduh|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
ItsThatGuyBrent|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
ItsThatGuyBrent|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
MomCat_Reviews|HillaryforOH|0.5983|0.103|0.665|0.232|"RT @HillaryforOH: Rose escaped Nazi Germany at 15 &amp; is a proud American! Despite a recent broken hip, she just proudly cast her ballot for"
JulieCTaylor|twitter|0.5859|0.0|0.833|0.167|Amazing that I never see reports of votes switching from Hillary to Trump. Always the other way. Makes me wonder.Hm https://t.co/yu85qCqIYp
justmyowndrama|Pamela_Moore13|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
justmyowndrama|twitter|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
Pick6_|s_tamikah|0.3182|0.0|0.905|0.095|"RT @s_tamikah: Men get a hold on these Women, cause Feminist gonna make sure Hillary win's JUST because she's not a Man&amp;if she doesn't the"
FLMENFORTRUMP|SonofLiberty357|0.4939|0.0|0.824|0.176|RT @SonofLiberty357: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/VpmqCeml3e
FLMENFORTRUMP|thegatewaypundit|0.4939|0.0|0.824|0.176|RT @SonofLiberty357: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/VpmqCeml3e
ty6939|DontTread_2nd|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
ty6939|twitter|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
LucasSchobert|CloydRivers|0.0|0.0|1.0|0.0|RT @CloydRivers: Hillary for President.Merica. https://t.co/PPkPj8mGEH
LucasSchobert|twitter|0.0|0.0|1.0|0.0|RT @CloydRivers: Hillary for President.Merica. https://t.co/PPkPj8mGEH
sfkaw69|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
MontriciaHubba1|wikileaks|-0.2732|0.139|0.861|0.0|RT @wikileaks: Its ignorant to vote for Hillary Clinton without reading WikiLeaks https://t.co/Tiywc9Nrgr https://t.co/c0QaJW4hCi
MontriciaHubba1|denverpost|-0.2732|0.139|0.861|0.0|RT @wikileaks: Its ignorant to vote for Hillary Clinton without reading WikiLeaks https://t.co/Tiywc9Nrgr https://t.co/c0QaJW4hCi
tlvrp_russia|therussophile|-0.2732|0.195|0.667|0.138|#Moscow #SaintPetersburg Stanford University Confirms Democratic 2016 Election Fraud In Favor of Hillary Clinton https://t.co/9Ps7WcZp6q
ttm2x|DJ_SKEME|0.7579|0.0|0.629|0.371|RT @DJ_SKEME: #BlackTwitter will be pure entertainment tonight whether Hillary or Trump wins
MayorSnart|Queentette|0.5996|0.069|0.701|0.23|@Queentette Hillary isn't a white straight male. So everything she does is ok. As long as she's not that scumbag Trump
xactnode|kincannon_show|-0.5849|0.296|0.704|0.0|RT @kincannon_show: This is very bad for Hillary --&gt; https://t.co/lv5ybXLiHZ
xactnode|twitter|-0.5849|0.296|0.704|0.0|RT @kincannon_show: This is very bad for Hillary --&gt; https://t.co/lv5ybXLiHZ
ViciousVeeeeeee|jozenc|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
ViciousVeeeeeee|twitter|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
jsirwin67|Stonewall_77|0.4847|0.0|0.851|0.149|"RT @Stonewall_77: If This Isn't Torture, What is?THIS is what Hillary Clinton explicitly defended at the third presidential debate."
doitlikeAmb|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Jennife40966102|USATODAY|0.4019|0.0|0.816|0.184|RT @USATODAY: Voters are pantsuit-ing up in support of Hillary Clinton. #ElectionNight https://t.co/puR0Ca8bbx
Jennife40966102|twitter|0.4019|0.0|0.816|0.184|RT @USATODAY: Voters are pantsuit-ing up in support of Hillary Clinton. #ElectionNight https://t.co/puR0Ca8bbx
arrowsmithwoman|WDFx2EU8|-0.3595|0.238|0.762|0.0|@WDFx2EU8 Bet there's no Hillary voters in that line!
kobybaker|TheOneandOnIyUS|0.7096|0.0|0.753|0.247|RT @TheOneandOnIyUS: The joke is on Hillary if she wins. She'll have to sit at the desk Monica sat under.
BULGEBULL|i2|0.4019|0.0|0.838|0.162|WATCH LIVE: Hillary Clinton and Donald Trump Hold Election Night Parties Only A Mile Apart  https://t.co/vGY5zOkGg6
viplive|tmz|0.0|0.0|1.0|0.0|Hillary and Donald -- Enough Already!!! You're Bleeding Us Dry https://t.co/5pXLd0oILP
DianaChavira6|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
DianaChavira6|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
beyoncedefense|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: .@Beyonce &amp;@S_C_ &amp;Hillary &amp;You?https://t.co/3TKJ4H68Kz https://t.co/DAxSZLuQUB
beyoncedefense|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: .@Beyonce &amp;@S_C_ &amp;Hillary &amp;You?https://t.co/3TKJ4H68Kz https://t.co/DAxSZLuQUB
karbob85|hardassettimes|0.5719|0.0|0.793|0.207|RT @hardassettimes: @BarbMuenchen @maggiebeauchamp All those people are certainly not waiting in line to vote for Crooked Hillary. Pray for
OdellSZN|StephForMVP30|0.7955|0.0|0.718|0.282|RT @StephForMVP30: If Trump or Hillary wins the election I'm moving out the country! Goodbye America and hello United States!
_khaliyaaah|AfroGumOfficiaI|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
_khaliyaaah|twitter|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
m_shepherd3|emilyo427|0.0|0.0|1.0|0.0|"RT @emilyo427: Same age, same stage of development, but only one has the right to life...makes sense right Hillary? https://t.co/FD35xt72wb"
m_shepherd3|twitter|0.0|0.0|1.0|0.0|"RT @emilyo427: Same age, same stage of development, but only one has the right to life...makes sense right Hillary? https://t.co/FD35xt72wb"
PastorTeeTalley|wiselatinaslink|0.4019|0.0|0.863|0.137|RT @wiselatinaslink: Hillary Clinton will treat women as equals. You know what Trump thinks of us. #ElectionNight https://t.co/jgMQt6sGbk
PastorTeeTalley|twitter|0.4019|0.0|0.863|0.137|RT @wiselatinaslink: Hillary Clinton will treat women as equals. You know what Trump thinks of us. #ElectionNight https://t.co/jgMQt6sGbk
GMWhiteAmerica|OnlineMagazin|-0.5267|0.207|0.714|0.079|RT @OnlineMagazin:  That made my day. Crooked Hillary supporter went into the trap when he wanted to steal the #DonaldTrump shield. ht
_Proud_American|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
thesessionista|AmberinSEA|0.9036|0.0|0.63|0.37|"@AmberinSEA I was thinking of you a few days ago, I remember how super pro-Hillary you were in 2008 at Genie!! Yay! (well, hopefully Yay!)"
dankpaul|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
dankpaul|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
AliceCoven|ChooseToBFree|-0.7506|0.39|0.61|0.0|"RT @ChooseToBFree: @ezinder Aiding and abetting the enemy IS treason, Sir. @HlLLARYCLINT0N#HillaryIndictment#HillarysEmails#Hillary#Dra"
Jaraselmanlol|JackJ|0.0772|0.0|0.894|0.106|@JackJ excuse me Hillary isn't any better... I'm out either way. #RIPAmerica
dahp0928|SoCal4Trump|0.0|0.0|1.0|0.0|"RT @SoCal4Trump: Bernie held a rally for Hillary today, but the student introducer went off script, trashed Hillary, and was led off stage."
Hacker_4_chan|LeighPatrick|0.0|0.0|1.0|0.0|"RT @LeighPatrick: Given the reports flooding in nationwide, you either vote Hillary or the machine votes Hillary for you. #Corruption #elec"
force4truth|ppetrov5|0.0|0.0|1.0|0.0|"RT @ppetrov5: Hillary Clinton and her campaign met with prioritiesUSA, which is against the law. #PodestaEmails35 #wikileaks #fbi https://t"
force4truth||0.0|0.0|1.0|0.0|"RT @ppetrov5: Hillary Clinton and her campaign met with prioritiesUSA, which is against the law. #PodestaEmails35 #wikileaks #fbi https://t"
debbiedo58|Nascar_Tom|-0.1111|0.148|0.719|0.133|RT @Nascar_Tom: STUPID pundit so called reporters really think If #CHEATINGHILLARY wins that WE THE PEOPLE HAVE to come together with Hilla
SweetFreedom29|CounterMoonbat|0.2023|0.128|0.677|0.195|RT @CounterMoonbat: Hillary smeared women who were assaulted and takes millions from regimes that treat women like property. Spare me the f
badmem_x86|Scarlett210|-0.765|0.28|0.72|0.0|"RT @Scarlett210: And #Hillary is a self-serving #elitist who'll continue #globalist policies, destroy ur safety&amp; deprive ur kids of a futur"
GraceRogerson_|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
GraceRogerson_|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
tkrobinson_|cjlake|-0.7506|0.381|0.619|0.0|RT @cjlake: I swear if FLOTUS doesn't pull a Hillary in a few terms...I'll cry. Fr. I'll cry.
JrmezaMeza|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
JrmezaMeza|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
JacksonJoshua73|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
JacksonJoshua73|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
humaneffect|twitter|-0.3595|0.185|0.815|0.0|Hillary NEEDS YOUR VOTE.Trump is getting Indiana.send a message now. no trump! https://t.co/dy4nAUJB06
amberhearrds||0.5267|0.0|0.761|0.239|can my early birthday present be Hillary Clinton as President please @ god @ the entire fucking country
rakiichak|officialSmith_|0.3612|0.0|0.783|0.217|RT @officialSmith_: *casts vote for Hillary*Hillary: Thank you s--Me: https://t.co/rmDqKBTo1i
rakiichak|twitter|0.3612|0.0|0.783|0.217|RT @officialSmith_: *casts vote for Hillary*Hillary: Thank you s--Me: https://t.co/rmDqKBTo1i
mvrleysky|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
mvrleysky|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
iamBoozforeal|rudeboyy|0.0772|0.0|0.902|0.098|Video: Common Freestyles About Hillary Clinton &amp; Voting On Election Day  https://t.co/GKLwSuEZI8 https://t.co/3vdRtLdzD4
erlckachaa|ConstanceQueen8|0.0|0.0|1.0|0.0|RT @ConstanceQueen8: Tracking Voter TurnOutHope This TrendsIn The Other 44 States#Vote4Trump #Defeat_Hillary#HillaryForPrisi
mykaela_watkins|Avstvn|-0.1695|0.196|0.804|0.0|"RT @Avstvn: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
iceman120|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
iceman120|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
elinepomstra|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
MooreAnthony12|TheWorldOfFunny|0.0|0.0|1.0|0.0|RT @TheWorldOfFunny: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/rYVq0sC4U5
MooreAnthony12|twitter|0.0|0.0|1.0|0.0|RT @TheWorldOfFunny: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/rYVq0sC4U5
itsbeenlit|NathanZed|0.5267|0.0|0.848|0.152|RT @NathanZed: my 7 year old cousin just now: is Hellen Keller winning me: whatcousin: Hellen Kellerme: Hillary Clinton? cousin: I dont
darylrjho|joshpan|0.0|0.0|1.0|0.0|RT @joshpan: what if i am hillary clinton
armadillobee|PrisonPlanet|0.4404|0.0|0.884|0.116|RT @PrisonPlanet: Hey Hillary supporters; You're about to vote for someone who is funded by countries that still execute gay people. How pr
Maddie_Mae4|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Maddie_Mae4|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
YewtreeGirl|rorysutherland|-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
YewtreeGirl||-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
Chrisspero1|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Chrisspero1|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
FortuneClint|youtube|0.0|0.0|1.0|0.0|Voting machines in Pennsylvania switch Trump votes to Hillary https://t.co/MB4HMHDGbb
robert_burrito|TheSometimesWhy|-0.7792|0.299|0.701|0.0|"@TheSometimesWhy but I know allowing Hillary is far worse. And if we don't agree, it is what it is"
tweetheart96_|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
tweetheart96_|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
DeplorableRich|TRay1949|0.0|0.0|1.0|0.0|RT @TRay1949: Hillary's Kissin KKK  https://t.co/2RoehKOfht
DeplorableRich|twitter|0.0|0.0|1.0|0.0|RT @TRay1949: Hillary's Kissin KKK  https://t.co/2RoehKOfht
amigoalfil|HillaryClinton|0.0772|0.0|0.942|0.058|"RT @HillaryClinton: ""Its not just my name or Donald Trumps name on the ballotits the kind of country we want. Hillary https://t.co/jf"
amigoalfil|t|0.0772|0.0|0.942|0.058|"RT @HillaryClinton: ""Its not just my name or Donald Trumps name on the ballotits the kind of country we want. Hillary https://t.co/jf"
CharlieEricks10|LarryT1940|0.0|0.0|1.0|0.0|RT @LarryT1940: #Vote4Trump and don't let these #Slime_balls of #Hillary's drive you away from voting. Your vote may push #Trump over the t
ReynoldHawthor2|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
GLuviano|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
nemyheartsmanga|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
nancy73gg|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
diaaanuuuh|SportsTakeJames|-0.1531|0.117|0.789|0.094|RT @SportsTakeJames: Choosing between Hillary &amp; Trump to replace Obama is like when the McDonald's ice cream machine is broken &amp; you gotta
juliann23_|elias_chairez|-0.2348|0.212|0.635|0.153|RT @elias_chairez: People giving Hillary their vote so Trump won't win: https://t.co/0SfLCKj03a
juliann23_|twitter|-0.2348|0.212|0.635|0.153|RT @elias_chairez: People giving Hillary their vote so Trump won't win: https://t.co/0SfLCKj03a
Julian_A_Cox|DESlRABLE|0.3453|0.078|0.779|0.143|@DESlRABLE @Calum5SOS Ya think that's weird? The other guy (Hillary's client) fancies himself as GOD! Get this athe https://t.co/rqIhMjbZH7
Julian_A_Cox|twitter|0.3453|0.078|0.779|0.143|@DESlRABLE @Calum5SOS Ya think that's weird? The other guy (Hillary's client) fancies himself as GOD! Get this athe https://t.co/rqIhMjbZH7
SprockDaddy|itsbillertime1|-0.6808|0.318|0.682|0.0|"RT @itsbillertime1: Donna Brazile cheats for Hillary, lies about it on live TV. https://t.co/6n94zv2bbP"
SprockDaddy|twitter|-0.6808|0.318|0.682|0.0|"RT @itsbillertime1: Donna Brazile cheats for Hillary, lies about it on live TV. https://t.co/6n94zv2bbP"
mcphersonfamily|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: Remember, Hillary is 46,000 votes behind Obama in just Pinellas County."
CollinsDionte|twitter|0.0|0.0|1.0|0.0|Hillary will still become POTUS regardless. https://t.co/zgyZkCTHg2
Kathywa48814788|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
Kathywa48814788|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
Jessicamertz4|RepCoriFournier|0.4404|0.0|0.879|0.121|RT @RepCoriFournier: Hmm... odd.... @CNN claims LATINOS are flooding the polls for Hillary. Funny how very diff LATINOS claim they feel abo
pllilje1|OnlineMagazin|-0.5267|0.207|0.714|0.079|RT @OnlineMagazin:  That made my day. Crooked Hillary supporter went into the trap when he wanted to steal the #DonaldTrump shield. ht
middlewingJeff|ClubBayern|-0.6369|0.345|0.5|0.155|RT @ClubBayern: Justice Poll: What's Hillary's worst crime? #ElectionDay #ElectionNight #WTFAmericaIn5Words #VotingDaySongs #MAGA #ivoted
leannelovsin|voguemagazine|0.0|0.0|1.0|0.0|"RT @voguemagazine: ""She doesnt realize it yet, but Election Day is a moment in history for both of us."" https://t.co/aP0pq0q274"
leannelovsin|vogue|0.0|0.0|1.0|0.0|"RT @voguemagazine: ""She doesnt realize it yet, but Election Day is a moment in history for both of us."" https://t.co/aP0pq0q274"
KeswickPinhead|SenFallon2016|0.2481|0.089|0.786|0.125|"RT @SenFallon2016: This election is rigged! I intended to vote for #Trump today, when Jesus smacked me upside the head &amp; made my hand vote"
ifollowcoby|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
ifollowcoby|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
xmoshingbatmanx|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
xmoshingbatmanx|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
xDrakeFam|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
xDrakeFam|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Chrisrlamar|DTorday|-0.4497|0.235|0.624|0.141|"@DTorday @JamesOKeefeIII @daveweigel but you're cheating the election for Hillary, so how is that fair?"
teenagefur|FlawlessDog|0.0|0.0|1.0|0.0|"RT @FlawlessDog: If you're in line before polls close, you have the right to vote. Stay in line and vote for Hillary. #ImWithHer"
hibadjedaini|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
henderson_mark|TurtleBoySports|0.7178|0.0|0.5|0.5|"@TurtleBoySports Wow, more surprised by early than Hillary."
jmhpa|RepCoriFournier|0.0|0.0|1.0|0.0|RT @RepCoriFournier: This is what @CNN is counting on with the BIG push on their network that Republicans will be voting HILLARY n republic
Worped4|ILoveBernie1|-0.8689|0.329|0.671|0.0|"RT @ILoveBernie1: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, https"
toddhenderson23|WayneDupreeShow|-0.296|0.136|0.864|0.0|RT @WayneDupreeShow:  Huckabee: Hillary Has No Empathy For The Working Class https://t.co/NEEjhHx6Zy #DrainTheSwamp #TrumpTrain https://t.
toddhenderson23|newsninja2012|-0.296|0.136|0.864|0.0|RT @WayneDupreeShow:  Huckabee: Hillary Has No Empathy For The Working Class https://t.co/NEEjhHx6Zy #DrainTheSwamp #TrumpTrain https://t.
KatEdmiston|BruceBartlett|0.6311|0.076|0.688|0.235|"RT @BruceBartlett: For the record, I voted enthusiastically for Hillary Clinton today. She may not be perfect, but she's light years better"
ChiefCRX340|BlastingNews|0.0|0.0|1.0|0.0|RT @BlastingNews: #election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR http
ChiefCRX340|us|0.0|0.0|1.0|0.0|RT @BlastingNews: #election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR http
DawnieRotten|worldnetdaily|0.4588|0.159|0.53|0.311|Hillary puts nation at great risk https://t.co/1FjeguvPjc via @worldnetdaily
DawnieRotten|wnd|0.4588|0.159|0.53|0.311|Hillary puts nation at great risk https://t.co/1FjeguvPjc via @worldnetdaily
tinymyg|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
guadss_|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
soleileva31|stephstabile8|0.0|0.0|1.0|0.0|RT @stephstabile8: trump &gt; hillary
chrisldoster|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
franco_dimuro|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
franco_dimuro|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
GBabySanch|twitter|0.0|0.0|1.0|0.0|My prediction: Hillary gonna put up numbers https://t.co/aQd3PgJw4E
WaltyAlvarez|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
miracles3337|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
miracles3337||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
steve62269|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
Filterlbc|AltStreamMedia|0.0258|0.139|0.717|0.143|"RT @AltStreamMedia: Judge to Trump: ""Only you can bring Hillary to justice. Our corrupt judicial system has failed, #LockHerUp"""
INFOS_EN|belfasttelegraph|0.25|0.0|0.824|0.176|US election results: Donald Trump and Hillary Clinton await their verdict of voters - Belfast Telegraph https://t.co/ypMwah7jqC
12aptor|kgarrison|-0.6876|0.296|0.582|0.122|RT @kgarrison: Republicans may be RINOS or weak kneed but they are not criminals like the Democrats. Democrats are dishonest which is why t
ekujpg|jacksfilms|0.0|0.0|1.0|0.0|RT @jacksfilms: You only have a few hours left to write your Trump/Hillary fanfiction
karbripal3|yankeebrit77|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
karbripal3|twitter|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
jwl868|BBCScotlandNews|0.0|0.0|1.0|0.0|RT @BBCScotlandNews: Holyrood leaders back Hillary Clinton for US president as the race for the White House draws to a close https://t.co/6
jwl868|twitter|0.0|0.0|1.0|0.0|RT @BBCScotlandNews: Holyrood leaders back Hillary Clinton for US president as the race for the White House draws to a close https://t.co/6
azakharov82|foreignpolicy|0.0|0.0|1.0|0.0|What Kind of President Will Hillary Clinton Be? | Foreign Policy https://t.co/mWXlnD4RrY
dwzd|HillaryClinton|0.0|0.0|1.0|0.0|@HillaryClinton I voted for Hillary ..Team Hillary!!!
_PinkkMoscato|beyupdates_|0.3612|0.0|0.815|0.185|RT @beyupdates_: Me: *votes for Hillary* Hillary: Thank you for vot-Me: https://t.co/nx99GlD5gc
_PinkkMoscato|twitter|0.3612|0.0|0.815|0.185|RT @beyupdates_: Me: *votes for Hillary* Hillary: Thank you for vot-Me: https://t.co/nx99GlD5gc
increase32|TravisRuger|-0.2263|0.203|0.642|0.155|RT @TravisRuger: A vote for Hillary is supporting election fraud.    #PodestaEmails33 #ElectionFinalThoughts #DNCLeaks2 #NeverHillary https
FlySince91_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
FlySince91_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ICollectCans|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
audreytan|FT|0.0|0.0|1.0|0.0|"RT @FT: As results come in, the polls point to a Hillary Clinton lead, but the race remains close in crucial swing states https://t.co/EQ1Q"
audreytan|t|0.0|0.0|1.0|0.0|"RT @FT: As results come in, the polls point to a Hillary Clinton lead, but the race remains close in crucial swing states https://t.co/EQ1Q"
hanxine|localblactivist|0.0|0.0|1.0|0.0|RT @localblactivist: Hillarys wrongdoings have gone unaccounted for in many instances. (ex. Clinton has been much more than a bit player i
MCGA2019|eagoodlife|-0.8748|0.625|0.375|0.0|@eagoodlife Hillary threatening to attack Russia? More scary https://t.co/bpTwnAZWI8
MCGA2019|twitter|-0.8748|0.625|0.375|0.0|@eagoodlife Hillary threatening to attack Russia? More scary https://t.co/bpTwnAZWI8
Hunter_Ash23|Pamela_Moore13|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
Hunter_Ash23|twitter|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
fvckmefenty|hosthetic|0.5945|0.0|0.812|0.188|"RT @hosthetic: Beyonc, Jay Z, Katy Perry, Lady Gaga and so many other huge celebrities have supported Hillary and Donald still has a chanc"
natalierose3123|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
natalierose3123|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
Liee4Trump|halsteadg048|0.0|0.0|1.0|0.0|"RT @halsteadg048: Hillary Clinton and her campaign met with prioritiesUSA, which is against the law. #PodestaEmails35 #wikileaks #fbi https"
CKlein5852|AdamsFlaFan|0.0|0.0|1.0|0.0|RT @AdamsFlaFan: Hillary Clinton Is Trouncing Trump With Her Ground Game According To Exit Poll via @politicususa https://t.co/Fa8OqrLYog
CKlein5852|politicususa|0.0|0.0|1.0|0.0|RT @AdamsFlaFan: Hillary Clinton Is Trouncing Trump With Her Ground Game According To Exit Poll via @politicususa https://t.co/Fa8OqrLYog
TayNicoole|WesVengeance7|0.296|0.0|0.891|0.109|RT @WesVengeance7: The joke is on Hillary if she wins.She'll have to sit at the desk Monica sat under.
sophia_bonoma|BruhhhComedy|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
sophia_bonoma|twitter|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
ChuckCollier76|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @MaddieAndMichi @enjoynChi @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE
babycats29|activist360|0.0|0.0|1.0|0.0|RT @activist360: Michael Moore is spot-on about all the reasons to vote for Hillary Clinton: She is going to make an incredible president.
imA_Creator|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
osu922|ChaseBurcher|-0.3612|0.122|0.878|0.0|"@ChaseBurcher I wouldn't put anything past Hillary. She already rigged the primary for herself, which the process started years ago"
KarolineMarquis|BruhhhComedy|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
KarolineMarquis|twitter|0.5719|0.0|0.748|0.252|RT @BruhhhComedy: Left = Me if Trump winsRight = Me if Hillary wins https://t.co/zJgSN9LpkW
RonaldMRivera|Boogie2988|-0.4019|0.172|0.828|0.0|RT @Boogie2988: Donald trump and Hillary clinton are both in a plane crash.  Who survives?....america.
AlexWeis3|twitter|0.0|0.0|1.0|0.0|If you are voting for Hillary the voting has changed. Its now tomorrow Rt to spread the word!!! https://t.co/C1JyMEsDP2
Juzwik|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Juzwik|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
rjber15|CTU279|0.6588|0.0|0.812|0.188|RT @CTU279: Great CTU volunteers out early this morning at Joseph Gallagher for Issue 108 and Hillary! @mcropper1 @EricGordon_CEO @ShariOB
asssophieyoung|NathanZed|0.5267|0.0|0.848|0.152|RT @NathanZed: my 7 year old cousin just now: is Hellen Keller winning me: whatcousin: Hellen Kellerme: Hillary Clinton? cousin: I dont
jason8a99|TheFunnyVine|0.0|0.0|1.0|0.0|RT @TheFunnyVine: Hillary out here trying to get the black vote https://t.co/x6lSCVIeGM
jason8a99|vine|0.0|0.0|1.0|0.0|RT @TheFunnyVine: Hillary out here trying to get the black vote https://t.co/x6lSCVIeGM
goawayitsnotme|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
DTharp1988|FoxNews|0.0|0.0|1.0|0.0|@FoxNews Some will vote for Hillary. Some will vote for Trump. Some will vote AGAINST Hillary or against Trump. I voted for my son's future.
theycallmegin|FemaleTexts|0.0|0.0|1.0|0.0|RT @FemaleTexts: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/Y01V5X3Als
theycallmegin|twitter|0.0|0.0|1.0|0.0|RT @FemaleTexts: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/Y01V5X3Als
Shhhh116|weknowwhatsbest|0.5574|0.097|0.672|0.231|"RT @weknowwhatsbest: Go easy on Hillary.  C'mon, be honest, I think we've all lied for 30 years at one time or another."
Michelle3wits|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
Michelle3wits|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
an_gonzalez22|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
yungjenz|NathanZed|0.5267|0.0|0.848|0.152|RT @NathanZed: my 7 year old cousin just now: is Hellen Keller winning me: whatcousin: Hellen Kellerme: Hillary Clinton? cousin: I dont
nrsbrnsff|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
nrsbrnsff|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
stticck|NeilTurner_|-0.6514|0.265|0.735|0.0|RT @NeilTurner_: @realDonaldTrump WE CAN PUT HILLARY IN PRISON BY VOTING TODAY! https://t.co/xSiV7G0kHQ
stticck|twitter|-0.6514|0.265|0.735|0.0|RT @NeilTurner_: @realDonaldTrump WE CAN PUT HILLARY IN PRISON BY VOTING TODAY! https://t.co/xSiV7G0kHQ
rcbbstcrk|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
Polysexuals|arzE|0.7865|0.0|0.729|0.271|RT @arzE: voting for Hillary doesn't have to be ur longest yeah boy ever. It can be ur shorter yeah boy ever. Just uhh don't waste ur yeah
lacey2123|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
lacey2123|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
sorryimspencerr|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Baskin_97|6PAPl|0.4404|0.0|0.879|0.121|RT @6PAPl: if kodak black believes hillary can do a good job with our country then we gotta go vote for hillary https://t.co/RWmwK8wHUR
Baskin_97|twitter|0.4404|0.0|0.879|0.121|RT @6PAPl: if kodak black believes hillary can do a good job with our country then we gotta go vote for hillary https://t.co/RWmwK8wHUR
Meghang622|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Meghang622|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
P1ssed_K1d|AlghamdiLife|0.7269|0.0|0.681|0.319|"@AlghamdiLife You're right, thanks to Hillary funding them all. Coming to an end my friend."
xoC_Lianne|TomiLahren|0.4717|0.0|0.861|0.139|RT @TomiLahren: If you're not voting for Trump don't you dare bitch when we get Hillary. Real talk. #MAGA #ElectionDay
xGoldiLOCKx|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
xGoldiLOCKx|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
jazminxrod|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: Florida, its Election Day! Polls are open from 7am-7pm. Confirm your polling place now and go vote for Hillary! https:"
meghanhollowayy|chasemylovex|-0.3586|0.127|0.873|0.0|"RT @chasemylovex: no, Hillary is not the ""ideal candidate"" but we still gonna vote for her tho... and we'll deal with sis later, ya hear me"
Helena_Vasc|nick_steinmetz|0.0|0.0|1.0|0.0|RT @nick_steinmetz: Suddenly broward goes 100% for Hillary https://t.co/qQhzFNo7SL
Helena_Vasc|twitter|0.0|0.0|1.0|0.0|RT @nick_steinmetz: Suddenly broward goes 100% for Hillary https://t.co/qQhzFNo7SL
leamjavier_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
idklife348|ridevocals|-0.4588|0.146|0.778|0.075|"RT @ridevocals: WHY ARE PEOPLE VOTING TRUMP BECAUSE ""HILLARY IS A CRIMINAL"" WHEN THE FBI ALREADY CLEARED HER AND TRUMP IS GOING TO COURT FO"
INFOS_EN|bustle|0.4019|0.0|0.838|0.162|"""Pantsuit Nation"" Stories About Voting For Hillary Clinton Offer A Home Stretch Election Boost - Bustle https://t.co/XFy9b3f4WW"
JacekJasinski|NTXShopping|0.5859|0.0|0.833|0.167|RT @NTXShopping: Hillary Clinton has enough electoral votes to win the White House in final Fix map https://t.co/HK9GdUvOn3 #ImWithHer #Str
JacekJasinski|linkis|0.5859|0.0|0.833|0.167|RT @NTXShopping: Hillary Clinton has enough electoral votes to win the White House in final Fix map https://t.co/HK9GdUvOn3 #ImWithHer #Str
Ebbi_Ling|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Ebbi_Ling|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Eag1e0ne|MarkDice|-0.4738|0.118|0.882|0.0|RT @MarkDice: Do Hillary voters have to fill out their ballots in blood?  Vote for Trump and let's send that witch into retirement!! #Elect
Juan_Migg|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
Juan_Migg|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
andregreen0|CNN|0.6369|0.0|0.833|0.167|"RT @CNN: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/QurbNzL1BK"
andregreen0|cnn|0.6369|0.0|0.833|0.167|"RT @CNN: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/QurbNzL1BK"
NotcoolOToole|TheTrumpPuppet|0.0|0.0|1.0|0.0|"RT @TheTrumpPuppet: ""Hello Hillary. How are you doing?"" #Trump #TheTrumpPuppet #Election #ElectionDay https://t.co/iPeB6nFXbl"
NotcoolOToole|vine|0.0|0.0|1.0|0.0|"RT @TheTrumpPuppet: ""Hello Hillary. How are you doing?"" #Trump #TheTrumpPuppet #Election #ElectionDay https://t.co/iPeB6nFXbl"
veeemariee_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
veeemariee_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
shotgunfetus|brobert545|0.25|0.06|0.84|0.1|"RT @brobert545: #Gaga and #HillaryClinton is it me, or does Hillary look like a crazed rodent? It takes a lot to make Gaga pretty... https:"
scarredbushido|Grummz|0.8689|0.078|0.523|0.399|@Grummz if hillary wins im avoiding watch TV because they keep going on about her being first female lol like i care.
Refinery29|refinery29|0.4588|0.0|0.75|0.25|How your favorite celebs are voting during #ElectionDay: https://t.co/OWRZ0dyO0m https://t.co/OyC6vTclZ9
confusednyy|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
confusednyy|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
babydulce_maria|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
babydulce_maria|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
brodyb_17|BasebalIy|0.0|0.0|1.0|0.0|RT @BasebalIy: Hillary bunts
jadedswine|twitter|0.0|0.0|1.0|0.0|Hillary Clinton = unaccomplished to the power of 30.https://t.co/0VLlxxnsmP #draintheswamp https://t.co/Wvc2G2ik8v
CariThumel|kylegriffin1|0.6369|0.0|0.846|0.154|"RT @kylegriffin1: Clinton camp out w/ new behind-the-scenes vids of HRC, best may be Bill jumping up and down after the 1st debate: https:/"
CariThumel||0.6369|0.0|0.846|0.154|"RT @kylegriffin1: Clinton camp out w/ new behind-the-scenes vids of HRC, best may be Bill jumping up and down after the 1st debate: https:/"
couchycraig|MagicRoyalty|0.3252|0.059|0.818|0.123|"RT @MagicRoyalty: Hillary doesn't want to #MAGA -- This makes Pepe sad.Please don't make Pepe sad, vote Trump.#ElectionDay https://t.c"
couchycraig||0.3252|0.059|0.818|0.123|"RT @MagicRoyalty: Hillary doesn't want to #MAGA -- This makes Pepe sad.Please don't make Pepe sad, vote Trump.#ElectionDay https://t.c"
KylarMartin|twitter|0.0|0.0|1.0|0.0|Would rather have Wild Bill from the Green Mile in office than Hillary. https://t.co/ItfJfnPJvk
AbbyMartinM|endingthefed|0.0|0.0|1.0|0.0|"WATCH  First Podesta Linked to SATANIC Rituals, Now THIS Breaks About Hillary! https://t.co/fHHEqkFE51 https://t.co/AfxWFGlTb3"
robertlesliejr|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
orBUMadBro|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
klarolinebonkai|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
klarolinebonkai|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Miss_Shanae_|lynnyChap|0.3887|0.0|0.893|0.107|"RT @lynnyChap: casted my ballot for Hillary and friends on Friday but if you haven't already, today is the day! VOTE VOTE VOTE! "
TengennToppa|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
TengennToppa|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
SlavichMadi|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
SlavichMadi|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
rosetaddie|LaziestCanine|-0.1695|0.196|0.804|0.0|"RT @LaziestCanine: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
valkgyria|sassytbh|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
valkgyria|twitter|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
DeathManagement|DrMartyFox|-0.296|0.121|0.879|0.0|RT @DrMartyFox: #ImVotingBecause We Must Stop DUAL #JUSTICEWhere #Deplorables Must Follow The #RuleOfLawWhile #Hillary &amp; Her Cronies
alexperns|iduitmann|0.5719|0.0|0.821|0.179|RT @iduitmann: joke's on Hillary if she wins. she'll have to sit at the desk Monica sat under.
racfink47|jamessmurray|0.3802|0.08|0.747|0.172|Screw Donald Trump and Hillary Clinton! @jamessmurray definitely has my vote cuz I believe in him
Mathiasian|SLandinSoCal|0.0|0.0|1.0|0.0|RT @SLandinSoCal: Does #Hillary have #Kuru? Contracted through #Canabalism. Symptoms mimic #Parkinsons. Would explain her inappropriate out
splash851851|JaredWyand|-0.7351|0.267|0.733|0.0|"RT @JaredWyand: WIKILEAKS RECAP#ImVotingBecause Hillary can't be allowed to lie, steal, &amp; cheat her way into the White House#ElectionFi"
stantheman3|YouTube|0.4084|0.0|0.767|0.233|VOTING AGAINST SATAN WORSHIPING HILLARY CLINTON 11/08/2016 https://t.co/5Z05hVYq5L via @YouTube
stantheman3|youtube|0.4084|0.0|0.767|0.233|VOTING AGAINST SATAN WORSHIPING HILLARY CLINTON 11/08/2016 https://t.co/5Z05hVYq5L via @YouTube
piercebboop|TheDonaldNews|0.627|0.0|0.708|0.292|RT @TheDonaldNews: LOOK AT CURRENT POPULAR VOTE!! TRUMP ==&gt;&gt; 6600  HILLARY===&gt;2043
MargaretMcgui16|worldnetdaily|0.516|0.0|0.836|0.164|"RT @worldnetdaily: CHURCH TAKES BOLD, ANTI-HILLARY STANCEPastor willing to give anyone a ride to polls, irrespective of vote https://t.co"
MargaretMcgui16|t|0.516|0.0|0.836|0.164|"RT @worldnetdaily: CHURCH TAKES BOLD, ANTI-HILLARY STANCEPastor willing to give anyone a ride to polls, irrespective of vote https://t.co"
reisegrrl1|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
Brisxyda|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
Brisxyda|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
haugherin|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
HanniaMorales1|twitter|-0.4939|0.222|0.696|0.082|Hillary: im not doing itThem: How bad do you want those votes? https://t.co/3lvQMPwvdW
NesUkijo|FalafelDad|-0.2617|0.089|0.911|0.0|RT @FalafelDad: When you can make billions by teaming up with Hillary but then you'd have to shake hands with a woman. https://t.co/O32PQPx
NesUkijo|t|-0.2617|0.089|0.911|0.0|RT @FalafelDad: When you can make billions by teaming up with Hillary but then you'd have to shake hands with a woman. https://t.co/O32PQPx
TheKidUnlifting|Saw_Insane|0.7579|0.0|0.667|0.333|RT @Saw_Insane: If Hillary Clinton wins I'm leaving America and going to the United States.
Ayethatsmera|CjayyTaughtHer|0.0|0.0|1.0|0.0|RT @CjayyTaughtHer: Trump Vs Hillary  https://t.co/e3XUMJbgFY
Ayethatsmera|twitter|0.0|0.0|1.0|0.0|RT @CjayyTaughtHer: Trump Vs Hillary  https://t.co/e3XUMJbgFY
DR_DRE_a|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
tlvrp_russia|therussophile|-0.5994|0.163|0.837|0.0|#Moscow #SaintPetersburg Jill Stein: we could slip into nuclear war in the blink of an eye if Hillary Clinton has  https://t.co/hfII9nUp2h
pithypisces|TeamTrump|0.7184|0.0|0.714|0.286|"RT @TeamTrump: Hillary only cares about power, money &amp; herself. @realDonaldTrump cares about YOU, the American people.https://t.co/vmaBF3"
NWONightmare|LatestAnonNews|0.0|0.0|1.0|0.0|"RT @LatestAnonNews: Hillary Clinton and her campaign met with @prioritiesUSA, which is against the law. #PodestaEmails34 https://t.co/B1Zfg"
NWONightmare|t|0.0|0.0|1.0|0.0|"RT @LatestAnonNews: Hillary Clinton and her campaign met with @prioritiesUSA, which is against the law. #PodestaEmails34 https://t.co/B1Zfg"
MiYeAmanda|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
Wilshe467711|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
DianeRainie1|farrightgregy|-0.6523|0.186|0.814|0.0|RT @farrightgregy: RT PhillyGOP: UPDATE: Ward 37-9 (North Philly): Poll workers handing out Hillary Lit INSIDE polling station. ILLEGAL #Vo
Razionnn|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
DeloresVallot|aduanebrown|0.0258|0.1|0.795|0.105|"RT @aduanebrown: Democrats are going crazy. Hillary was supposed to shatter the glass ceiling tonight, looks like Trumps shattering the Dem"
AdrianConradie|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
AdrianConradie|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
charles_tindol|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
angiekelly4|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
angiekelly4|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
Peraltafqw|ml|0.3182|0.134|0.63|0.236|Don't take life to seriously :) #nyvotes Hillary o Trump https://t.co/NTS4bGxIpA
phyllisinirmo|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
lantetrain|ImKateCrawford|0.8309|0.0|0.72|0.28|RT @ImKateCrawford: #ElectionNight #Election2016 to all my American peeps for the love of sweet baby J get out and vote for Hillary!! #ImWi
echoezofsilence|jaureologist|-0.0516|0.207|0.591|0.202|RT @jaureologist: I DON'T CARE HOW MUCH Y'ALL HATE BOTH CANDIDATES YOU WILL VOTE FOR HILLARY WHETHER YOU LIKE IT OR NOT I REFUSE TO LET TRU
BrianRodd6|RealPika|0.4926|0.0|0.79|0.21|RT @RealPika: Pikachu would be better than Donald Trump and Hillary Clinton! https://t.co/Q5ZdbSHID2
BrianRodd6|twitter|0.4926|0.0|0.79|0.21|RT @RealPika: Pikachu would be better than Donald Trump and Hillary Clinton! https://t.co/Q5ZdbSHID2
Samasterrr|marwannafuq|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
Samasterrr|twitter|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
KenValliere|scottkutach|0.0|0.0|1.0|0.0|"RT @scottkutach: BREAKING:  CNN has just called Mexico, Syria, Iran, Saudi Arabia, Qatar &amp; Morocco for Hillary. #ElectionDay #MyVote2016"
hmay26|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
hmay26|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
doodlebug2102|umpire43|-0.8286|0.327|0.673|0.0|RT @umpire43: Machines in all battleground states are flipping votes to Hillary. Some are using fraction counting fraud. DEMAND A PAPER BAL
hillwarner|sassytbh|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
hillwarner|twitter|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
debra_bonanno|Vote3Fortrump|0.4404|0.0|0.775|0.225|RT @Vote3Fortrump: Leftist Hillary Supporters TOTALLY TRASHED Independence Hall https://t.co/V1rV5hXd9g https://t.co/ccVCGyDLYi
debra_bonanno|thefederalistpapers|0.4404|0.0|0.775|0.225|RT @Vote3Fortrump: Leftist Hillary Supporters TOTALLY TRASHED Independence Hall https://t.co/V1rV5hXd9g https://t.co/ccVCGyDLYi
TheGiantHogweed|clmazin|-0.8442|0.302|0.698|0.0|"RT @clmazin: ""Fail Bigly"" (2031) - Barry Pepper stars as failed Republican nominee Donald J. Trump in the story of his historic loss to Hil"
MostLikelyCunt|TheRealistMi|-0.6596|0.265|0.675|0.06|RT @TheRealistMi: Ppl died for you dumb ass ignorant ppl to vote and y'all keep saying how your not  Yea Hillary a liar but so are you.
shanda4real|ELLEmagazine|0.0|0.0|1.0|0.0|"RT @ELLEmagazine: Rihanna #ElectionDay outfit is everything, of course: https://t.co/nmAzf43qlb"
shanda4real|elle|0.0|0.0|1.0|0.0|"RT @ELLEmagazine: Rihanna #ElectionDay outfit is everything, of course: https://t.co/nmAzf43qlb"
Ky_serna5257|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Ky_serna5257|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
YOCUMILA|chanddlerriggs|0.0|0.0|1.0|0.0|RT @chanddlerriggs: boys at my school: feminists are so triggered over everything lolme: i would rather have hillary than trumpboys at
BlazinHope|StarbucksSanae|0.2146|0.378|0.291|0.33|"@StarbucksSanae NO, DON'T LET TRUMP WIN, NO, DON'T LET HILLARY WIN! WE'RE SCREWED!"
FashBoyHeyGirl|refinery29|0.0|0.0|1.0|0.0|Rihanna Has A Message For All You Non-Voters https://t.co/XieHxg0ASm
casey____bug|twitter|0.5994|0.0|0.62|0.38|Oh my god people at me work likes hillary..fuck https://t.co/Mfyfqe74Zd
Moviewatcher21|worldnetdaily|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
Moviewatcher21|wnd|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
Givenchy_beauty|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
Givenchy_beauty|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
RhiannonN14|pantsuitnation|0.7088|0.0|0.671|0.329|RT @pantsuitnation: Hillary Clinton thanks #pantsuitnation for our support! #werewithher #sheswithus https://t.co/o7Pu89jE8s via @thr
RhiannonN14|hollywoodreporter|0.7088|0.0|0.671|0.329|RT @pantsuitnation: Hillary Clinton thanks #pantsuitnation for our support! #werewithher #sheswithus https://t.co/o7Pu89jE8s via @thr
Kkowen400Keith|GMA|-0.1027|0.203|0.636|0.161|@GMA at gma your lack of objective reporting and trying to rig election with your hillary favored reports by the minute get ready to suck it
JcEmery9|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
JcEmery9|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
dcfriend3|twitter|0.0|0.0|1.0|0.0|Boohoo-wait until president Trump starts investigating Hillary and all the others mentioned in the #wikileaks relea https://t.co/sBjizsa0kZ
AlyviaHagearty|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
AlyviaHagearty|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
ilahi__|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
ilahi__|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
beth_macgill|arzE|0.7865|0.0|0.729|0.271|RT @arzE: voting for Hillary doesn't have to be ur longest yeah boy ever. It can be ur shorter yeah boy ever. Just uhh don't waste ur yeah
alpha_joe86|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
00LovelyDay00|vivelafra|0.0|0.0|1.0|0.0|RT @vivelafra: ATTENTION #TRUMPTRAIN: The MSM narrative is beginning to CRUMBLE.  States long given to #Hillary are now back in the toss-up
meganderson01|toriking68|0.7845|0.0|0.717|0.283|RT @toriking68: Everyone bashes Trump like Hillary is any better and everyone bashes Hillary like Trump is any better...in the end we're al
PMgeezer|LeighPatrick|0.0|0.0|1.0|0.0|"RT @LeighPatrick: Given the reports flooding in nationwide, you either vote Hillary or the machine votes Hillary for you. #Corruption #elec"
NoleTuff|POTUS|0.2023|0.0|0.921|0.079|@POTUS And on top of that while you're campaigning for Hillary all of America is paying for it with tax dollars.    Smfh
coolinit81|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
coolinit81|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
kennethmac2000|bbc|0.0|0.0|1.0|0.0|BBC News - Scottish leaders back Hillary Clinton for US president https://t.co/E6hW3SJ0lW
Philfandan|BocaRatonRC|0.4404|0.0|0.854|0.146|RT @BocaRatonRC: Who better to torch Hillary to a crisp on election eve than firebrand Tomi Lahren? https://t.co/rnfeyqgAOD https://t.co/4Z
Philfandan|bizpacreview|0.4404|0.0|0.854|0.146|RT @BocaRatonRC: Who better to torch Hillary to a crisp on election eve than firebrand Tomi Lahren? https://t.co/rnfeyqgAOD https://t.co/4Z
raymarin96|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
raymarin96|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ArianneCiana|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
gravenoise|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
tlvrp_russia|therussophile|0.0|0.0|1.0|0.0|#Moscow #SaintPetersburg Hillary Clinton: A Cabinet Full of Old World Nationalists and Information Operations In C https://t.co/lTgxBfCyzJ
lamaramironova4|cosmopolitan|0.0|0.0|1.0|0.0|Disability-Rights Activist Anastasia Somoza Casts Her Vote for Hillary Clinton https://t.co/r3sZFgLMEi https://t.co/wbjUdkzZyg
alex__dalton96|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
alex__dalton96|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
OliviaArntzen|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
DevanMcCormick|JeffersJordan|0.0772|0.0|0.925|0.075|RT @JeffersJordan: Knowing that people are actually voting for Hillary Clinton makes me want to throw up.
dylanulloaaa|OmniDestiny|0.1027|0.114|0.759|0.128|"RT @OmniDestiny: If Hillary wins and you're trying to get laid, there will probably be a lot of depressed Trumple chicks at the bars tonigh"
Xamerican|MariaYes2trump|0.81|0.108|0.514|0.378|RT @MariaYes2trump: TRUMP VOTER LINES ARE HUGE! THERE IS NO WAY HILLARY CAN LEGALLY WIN! https://t.co/ImNnufMQAi via @wordpressdotcom
Xamerican|themarshallreport|0.81|0.108|0.514|0.378|RT @MariaYes2trump: TRUMP VOTER LINES ARE HUGE! THERE IS NO WAY HILLARY CAN LEGALLY WIN! https://t.co/ImNnufMQAi via @wordpressdotcom
zeabraa|polaroidbones|-0.607|0.184|0.816|0.0|RT @polaroidbones: DONT SPLIT THE DEMOCRATIC VOTE TOMORROW CAUSE YOU DONT WANNA BE STUCK HILLARY OR TRUMP! ITS ONLY GONNA LEAVE US WITH TRU
_crystaalc|foreverjournie|0.7996|0.0|0.411|0.589|RT @foreverjournie: I really hope Hillary wins. #ElectionNight
maxxbadazzent|GLOGangHQ|0.0|0.0|1.0|0.0|RT @GLOGangHQ: Donald Trump Hillary Clinton Chief Keef GO VOTE TODAY CHIEF KEEF 4 PRESIDENT #Election2016 #MyVote2016 https://t.co/
maxxbadazzent|t|0.0|0.0|1.0|0.0|RT @GLOGangHQ: Donald Trump Hillary Clinton Chief Keef GO VOTE TODAY CHIEF KEEF 4 PRESIDENT #Election2016 #MyVote2016 https://t.co/
Chrissy06699126|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Chrissy06699126|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Lofdaproduction|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Lofdaproduction|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Mom74548299|ConstanceQueen8|0.0|0.0|1.0|0.0|RT @ConstanceQueen8: Tracking Voter TurnOutHope This TrendsIn The Other 44 States#Vote4Trump #Defeat_Hillary#HillaryForPrisi
peachymarz|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
selinakrieg|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
LostChicInPa|hermanbutler1|0.6369|0.0|0.729|0.271|"RT @hermanbutler1: The Miami Herald Endorses Hillary Clinton In A Simple, Yet Powerful Editorial https://t.co/fUFxhvPFhI #TNTweeters #USLat"
LostChicInPa|linkis|0.6369|0.0|0.729|0.271|"RT @hermanbutler1: The Miami Herald Endorses Hillary Clinton In A Simple, Yet Powerful Editorial https://t.co/fUFxhvPFhI #TNTweeters #USLat"
ra_estella|religiouscaviar|0.743|0.0|0.751|0.249|"RT @religiouscaviar: Hillary's been serving looks since the 60s, and tonight she'll serve Trump and his supporters by winning the presidenc"
calvalais|ProgtopiaBooks|0.0|0.0|1.0|0.0|RT @ProgtopiaBooks: Some Pittsburgh machines changing from Trump to Hillary.Problems call 1-866-OUR-VOTE
inafutureage|rorysutherland|-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
inafutureage||-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
Victoriaabeni|arzE|0.7865|0.0|0.729|0.271|RT @arzE: voting for Hillary doesn't have to be ur longest yeah boy ever. It can be ur shorter yeah boy ever. Just uhh don't waste ur yeah
Tommy_Reason|twitter|0.5719|0.0|0.654|0.346|Me if Trump wins:Me if Hillary wins: https://t.co/jbKJp1LaBw
notbapecamo|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
notbapecamo|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
sofiadaviddd|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
jennyy882|memeprovider|-0.1695|0.196|0.804|0.0|"RT @memeprovider: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
march4progress|rtyson82|-0.8883|0.451|0.549|0.0|RT @rtyson82: I'm mocking ALL crying Hillary supporters!Remember when you mocked Bernie delegates for crying at the convention?Karma 
larryqqueen|BradThor|0.4767|0.092|0.712|0.197|"RT @BradThor: I did not vote for the Orange Raccoon, nor did I vote for Corrupt Hillary Clinton. I voted Third Party and am damn proud of i"
P2017G|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
JulieMre|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
JulieMre|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
lovelyNovaBean|mitchellvii|0.5719|0.0|0.856|0.144|"RT @mitchellvii: Right now, Hillary is running roughly 60% behind Obama's performance in Hillsborough. Obama won FL in 2012 by only 1%. Dev"
livtompkins||-0.7603|0.266|0.734|0.0|"@ all my Redding followers, the Democratic tent apparently had a Hillary cutout wearing a Make America Nasty again shirt and I MISSED IT"
Danieljackson94|Michael_Goggans|0.0|0.0|1.0|0.0|RT @Michael_Goggans: All I know is if someone at my rank did what Hillary did they'd be in Leavenworth for 20+ years.
LuffyHS|FeaRMoho|0.0|0.0|1.0|0.0|@FeaRMoho i bet money that Hillary will not Receive 50% of the vote and i was offered 50% of my money that i bet.so i bet 1K i get 1.5K back
alinatede|tpolitical_news|-0.2263|0.112|0.888|0.0|RT @tpolitical_news: Navy veteran walks three blocks on crutches to vote for Hillary Clinton https://t.co/LyFduaFekQ https://t.co/pam7X1yIsu
alinatede|dailynewsbin|-0.2263|0.112|0.888|0.0|RT @tpolitical_news: Navy veteran walks three blocks on crutches to vote for Hillary Clinton https://t.co/LyFduaFekQ https://t.co/pam7X1yIsu
_Timone|ClarenceJWhite|0.0|0.069|0.863|0.069|RT @ClarenceJWhite: I feel like Trump &amp; Hillary are two divorced parents fighting over custody of us but we kinda just wanna go live with g
AlissaLeighh_|__ImNotReal__|0.1779|0.088|0.797|0.116|RT @__ImNotReal__: No we're voting against trump cause he's a despicable human being. If we had a better option than Hillary we'd vote agai
Indiiaaa15|polaroidbones|-0.607|0.184|0.816|0.0|RT @polaroidbones: DONT SPLIT THE DEMOCRATIC VOTE TOMORROW CAUSE YOU DONT WANNA BE STUCK HILLARY OR TRUMP! ITS ONLY GONNA LEAVE US WITH TRU
FacedHailz|SpeedKirbyX|0.3546|0.093|0.721|0.187|@SpeedKirbyX I think Hillary might be a great president because his husband didn't bring terrorist in America or start world war but he is a
kevhazel33|foxandfriends|0.5927|0.0|0.806|0.194|"RT @foxandfriends: .@GovMikeHuckabee: Hillary Clinton needs celebrities to get a crowd, but Donald Trump's supporters aren't coming for a f"
pacasandrs|realDonaldTrump|0.5574|0.0|0.816|0.184|@realDonaldTrump @BigDuhie1955 Vote Vote.Prove the MSM wrong.Every single vote counts.Hillary cannot change the balance of Supreme Court
YoungZlaw|_dbrand|0.0|0.0|1.0|0.0|RT @_dbrand: @cbaker92redskin @_willcompton Hillary wants to change our name
coldplayitcool|jaureologist|-0.0516|0.207|0.591|0.202|RT @jaureologist: I DON'T CARE HOW MUCH Y'ALL HATE BOTH CANDIDATES YOU WILL VOTE FOR HILLARY WHETHER YOU LIKE IT OR NOT I REFUSE TO LET TRU
tjhutson|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
tjhutson|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
RickAndKim30yrs|ReturnofRV|0.1779|0.109|0.746|0.144|"RT @ReturnofRV: Why are all the Hillary supporters, Hillary trolls, and Hillary mainstream media pundits strangely quiet?"
kiamarie30|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
MissLiberty1776|BoSnerdley|-0.4767|0.171|0.829|0.0|RT @BoSnerdley: WikiLeaks says it was under 'unrelenting' cyber attack on Election Day https://t.co/kf31Wxmlad via @MailOnline
MissLiberty1776|dailymail|-0.4767|0.171|0.829|0.0|RT @BoSnerdley: WikiLeaks says it was under 'unrelenting' cyber attack on Election Day https://t.co/kf31Wxmlad via @MailOnline
richeyyriann|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
richeyyriann|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
kristinaswaffo1|PriceParker2|-0.8126|0.346|0.654|0.0|"RT @PriceParker2: If voting for Trump makes you a racist, does voting for Hillary make you a criminal?"
jimveejr|prupaine|-0.7213|0.401|0.599|0.0|Vote to STOP HILLARY and an Incompetent GOP https://t.co/urRvFwscYH via @prupaine
jimveejr|prudencepaine|-0.7213|0.401|0.599|0.0|Vote to STOP HILLARY and an Incompetent GOP https://t.co/urRvFwscYH via @prupaine
illestclev|AweeBurrEee|-0.8594|0.263|0.737|0.0|RT @AweeBurrEee: people who oppose Hillary talk about her stance on abortion but won't discuss Trump's child rape case?????? babies are bab
throughthatmist|ilysmarigrande|0.6393|0.076|0.7|0.224|"RT @ilysmarigrande: Hillary might not be the best candidate, but u can't deny that she's better than Trump. I urge you to vote tomorrow. #I"
Toridevon|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
Toridevon|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
TJrasar|WaysThingsWork|0.1695|0.0|0.886|0.114|RT @WaysThingsWork: Obama endorsing Hillary and bashing trump? Let's not forget about this https://t.co/olDwdXaYFB
TJrasar|twitter|0.1695|0.0|0.886|0.114|RT @WaysThingsWork: Obama endorsing Hillary and bashing trump? Let's not forget about this https://t.co/olDwdXaYFB
tlvrp_russia|therussophile|-0.6908|0.322|0.678|0.0|"#Moscow #SaintPetersburg WikiLeaks criticizes both Hillary Clinton and Donald Trump, condemns McCarthyite Russia https://t.co/LWkUgemgl5"
beccaboiteau|CloydRivers|0.0|0.0|1.0|0.0|RT @CloydRivers: Im not against a woman bein President. Im just against that woman bein Hillary Clinton. Merica.
RadicalRW|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
leelamchop|LiberalLogic123|0.0|0.0|1.0|0.0|RT @LiberalLogic123: Reasons not to vote for Hillary:1. Chris Stevens2. Sean Smith3. Glen Doherty4. Tyrone Woods#ElectionFinalThough
_evaax0|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_evaax0|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
JessicainNYC|HillaryIn2016|0.0|0.0|1.0|0.0|RT @HillaryIn2016: My electoral vote predictionWinner: HillaryTime Race Will be Called: 8-8:15pmPTSenate: Dems WinHouse: GOP Wins#ImWi
_baileefox_|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
_baileefox_|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
HomerWhite|NewtTrump|-0.7269|0.316|0.575|0.109|RT @NewtTrump: RETWEET THIS LIKE CRAZY: Hillary's guilty of 70-100 violations of the US Constitution's Emoluments Clause and the media refu
meganmcginnis_|Awxme|-0.0387|0.057|0.943|0.0|RT @Awxme: Hillary Clinton may be the first f president. Sorry I meant to say female but the emale got deleted #ElectionDay
z1o9z6e9|NPR|0.0|0.0|1.0|0.0|RT @NPR: A spokesman for former President George W. Bush confirms to NPR that he and his wife voted for neither Donald Trump nor Hillary Cl
mlogika1|abcnews|0.25|0.0|0.867|0.133|RT @abcnews: .@HillaryClinton one step away from snaring her dream job #Election2016 https://t.co/XpMh9z93OP https://t.co/mPAFkHucrD
mlogika1|abc|0.25|0.0|0.867|0.133|RT @abcnews: .@HillaryClinton one step away from snaring her dream job #Election2016 https://t.co/XpMh9z93OP https://t.co/mPAFkHucrD
Hay_Bales23|EWT2015|-0.5106|0.268|0.732|0.0|RT @EWT2015: Hillary for prison 2016 #HillaryForPrison2016 #VeteransDay #vetslivesmatter #Election2016
GiselaHaaase|MANOUSHactress|-0.5423|0.127|0.873|0.0|RT @MANOUSHactress: if HILLARY will be president Germanys ANGELA MERKEL will be so deep up her ass that Hillary will be able to taste her @
JRayM5|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
JRayM5|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
kenzdelrey|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
itistj1|twitter|0.7865|0.0|0.565|0.435|What Hillary will look like when she realizes TRUMP WON  https://t.co/td3SM5IFgt
factanonverba7|marklevinshow|0.0|0.0|1.0|0.0|"RT @marklevinshow: Members of the jury, what do you say? https://t.co/mIRPiKFIWD"
factanonverba7|nationalreview|0.0|0.0|1.0|0.0|"RT @marklevinshow: Members of the jury, what do you say? https://t.co/mIRPiKFIWD"
tam_raww|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
tam_raww|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
oxnfre|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
LaneMorrow10|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
LaneMorrow10|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
eschwent|RobinDavani|-0.8941|0.339|0.661|0.0|RT @RobinDavani: @celestemc @CNNPolitics MORE VOTER FRAUD IN DURHAM COUNTY NC! 90 MINUTE EXTENSION TO CAST FRAUDULENT VOTES FOR HILLARY ALL
EnnisBruhh|DaiIyRap|0.0772|0.0|0.86|0.14|RT @DaiIyRap: Hillary Clinton doing the Mannequin Challenge https://t.co/yZXFZ1hNrn
EnnisBruhh|twitter|0.0772|0.0|0.86|0.14|RT @DaiIyRap: Hillary Clinton doing the Mannequin Challenge https://t.co/yZXFZ1hNrn
RobertD89815787|Scarlett210|-0.6597|0.234|0.766|0.0|RT @Scarlett210: If U can vote 4 #Hillary when you KNOW she's seriously ill maybe U shld forget ur enormous #Obamacare payt &amp; go to the hos
_arivna|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
ravensfan4|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
ravensfan4|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
katkrchniak|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
LKGNanci|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
Karaszewski|twitter|0.8126|0.0|0.72|0.28|If Hillary wins we are going to drink the Blue Label... if Trump wins we are going to drink everything https://t.co/t4Sr6HnCe1
TaraaTanner|Chubz3261|-0.5291|0.387|0.613|0.0|RT @Chubz3261: Hillary sucks but not like Monica #trumptrain
fuxkniaal|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
X5MSport15|Pamela_Moore13|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
X5MSport15|twitter|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
lulupink12|lois_rogers|0.8122|0.0|0.619|0.381|RT @lois_rogers: PHOTOS: #Hillary supporters trash lawn outside Independence Hall. They're so superior. https://t.co/ORs81FmXRO
lulupink12|theamericanmirror|0.8122|0.0|0.619|0.381|RT @lois_rogers: PHOTOS: #Hillary supporters trash lawn outside Independence Hall. They're so superior. https://t.co/ORs81FmXRO
timnemec|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
timnemec|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
_take_on_me_|CNN|0.0|0.0|1.0|0.0|RT @CNN: Watch 1993 footage of Bill and Hillary Clinton discussing the possibility of a woman running for president https://t.co/73tjhwsOUe
_take_on_me_|cnn|0.0|0.0|1.0|0.0|RT @CNN: Watch 1993 footage of Bill and Hillary Clinton discussing the possibility of a woman running for president https://t.co/73tjhwsOUe
MizCoretta|RedApplePol|0.5473|0.0|0.531|0.469|RT @RedApplePol: HERE'S HOPING  https://t.co/v0Yvnpt9hh
MizCoretta|aljazeera|0.5473|0.0|0.531|0.469|RT @RedApplePol: HERE'S HOPING  https://t.co/v0Yvnpt9hh
BenschoterKeith|lhfang|0.0|0.0|1.0|0.0|"RT @lhfang: Hillary watching the returns at a luxury hotel that costs up to $1,500 per night for a room https://t.co/vhlsFhYhbg"
BenschoterKeith|twitter|0.0|0.0|1.0|0.0|"RT @lhfang: Hillary watching the returns at a luxury hotel that costs up to $1,500 per night for a room https://t.co/vhlsFhYhbg"
KaisleXY|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
KaisleXY|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
hxrrera13|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
oxtilweoverdose|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
belladamaxx_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
hvilmary|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
hvilmary|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
LyndaJoHunt|jaynordlinger|0.7579|0.0|0.745|0.255|"RT @jaynordlinger: Hillary = luckiest politician ever. I know the hour is late, but are we SURE that Trump was not a Clinton plant?"
Suenorr11888815|FoxNews|0.0|0.0|1.0|0.0|RT @FoxNews: Crowds gathering for Hillary Clinton outside the Javits Center in New York City #ElectionNight #FoxNews2016 https://t.co/EdH4
Suenorr11888815|t|0.0|0.0|1.0|0.0|RT @FoxNews: Crowds gathering for Hillary Clinton outside the Javits Center in New York City #ElectionNight #FoxNews2016 https://t.co/EdH4
gabbie_4223|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
RM3Barcelona4|Chappynash|-0.6705|0.234|0.766|0.0|"RT @Chappynash: @SamWiseSW Hillary is worse.  She will flip the SCOTUS into a legislative judiciary for a generation. Trump is a jerk, she"
stairwaylover|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
stairwaylover|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
greenlawley|lovelaurenxjenn|0.5719|0.0|0.821|0.179|RT @lovelaurenxjenn: If Trump or Hillary  Wins The Election I Am Moving  Out Of The Country  Goodbye America  Hello   N
FilipDobi|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
peaceharmony16|Vets_Vs_Trump|0.7404|0.0|0.77|0.23|@Vets_Vs_Trump @PAMsLOvE @MorganLsneed YOU SURE CAN BREAK THE LAW AND GET AWAY FROM IT LIKE HILLARY . THAT IS WHAT YOU ARE GOING FOR
davidysteph|twitter|0.0|0.0|1.0|0.0|"6:59 in the VA suburbs, one minute before pools close. I just knocked on my last door canvassing for Hillary. Pleas https://t.co/ekOCYXuZgs"
RossGoldband|Redistrict|0.6908|0.0|0.778|0.222|"RT @Redistrict: Just one final thing: Remember, whatever the popular vote margin tonight, it should be ~1.5% better for Hillary Clinton by"
KaceyIlliot1669|jaketapper|-0.8687|0.376|0.542|0.081|"@jaketapper Trump is the only choice for us! Hillary cheats, lies and steals. She even cheated at the debates with help from CNN"
xohannah__|porn_horse|-0.7656|0.292|0.708|0.0|RT @porn_horse: Hillary campaigner employed FORBIDDEN MAGIC to do a kickflip in heels. No one is talking about this!!!https://t.co/GD9L0u
xohannah__|t|-0.7656|0.292|0.708|0.0|RT @porn_horse: Hillary campaigner employed FORBIDDEN MAGIC to do a kickflip in heels. No one is talking about this!!!https://t.co/GD9L0u
woIfbitch|JoshBasiliTV|-0.0516|0.224|0.51|0.265|@JoshBasiliTV please tell me u voted for hillary the devil its our only hope
trippyy__manee|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
mi4of5jaa|BruceBartlett|0.6311|0.076|0.688|0.235|"RT @BruceBartlett: For the record, I voted enthusiastically for Hillary Clinton today. She may not be perfect, but she's light years better"
Mrgee_bande|Ary_AntiPT|0.0|0.0|1.0|0.0|"RT @Ary_AntiPT: Trump up 70.5% to Hillary's 25.8% in Indiana. 35,646 votes to 13,049 #ElectionNight"
Kovach727|lizcgoodwin|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
Kovach727|twitter|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
roberpesca|FrankLuntz|0.6369|0.0|0.733|0.267|"RT @FrankLuntz: The numbers I'm getting now suggest a nationwide turnout that strongly favors Hillary.And if Hillary does well, so will d"
tiamomv|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
XicanoAdrian|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
XicanoAdrian|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
theOGericmullin|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
novelparadise|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
novelparadise|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Wbkirkendall|BlissTabitha|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
Wbkirkendall|weaselzippers|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
TheGwardian|OmniDestiny|0.1027|0.114|0.759|0.128|"RT @OmniDestiny: If Hillary wins and you're trying to get laid, there will probably be a lot of depressed Trumple chicks at the bars tonigh"
She_is_morg|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
She_is_morg|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
KailynnPerkins|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
KailynnPerkins|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Sxlcedo|TheBardockObama|0.4215|0.0|0.833|0.167|"RT @TheBardockObama: ""And your new president of the United States of America, Hillary Clinton""Hillary: https://t.co/9SPo9UJ6ig"
Sxlcedo|twitter|0.4215|0.0|0.833|0.167|"RT @TheBardockObama: ""And your new president of the United States of America, Hillary Clinton""Hillary: https://t.co/9SPo9UJ6ig"
Jennife51072808|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
my6girls2012|PrisonPlanet|-0.5563|0.204|0.796|0.0|RT @PrisonPlanet: #SpiritCooking turned out to be more damaging to Clinton than Comey's bluff. https://t.co/m4juc4F2dR
my6girls2012|thegatewaypundit|-0.5563|0.204|0.796|0.0|RT @PrisonPlanet: #SpiritCooking turned out to be more damaging to Clinton than Comey's bluff. https://t.co/m4juc4F2dR
plasmagender|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
E46lopez|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
E46lopez|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
creminsmom|MCrisCardena|-0.4003|0.119|0.881|0.0|@MCrisCardena If Hillary worked for a bank (any US Company) &amp;  released Confidential Info.... She is fired.... Fire Hillary .... Vote Trump!
NormandinRob|trump_florida|0.4019|0.0|0.828|0.172|RT @trump_florida: Source: The Military Times951 Active Duty Troops PolledTrump 54%     Hillary 25%#TrumpPence16 https://t.co/t1n374qx7M
NormandinRob|twitter|0.4019|0.0|0.828|0.172|RT @trump_florida: Source: The Military Times951 Active Duty Troops PolledTrump 54%     Hillary 25%#TrumpPence16 https://t.co/t1n374qx7M
amigoalfil|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: ""If you believe in science and that we have to act on climate change, then you have to vote!"" Hillary https://t.co/jfd"
amigoalfil|t|0.0|0.0|1.0|0.0|"RT @HillaryClinton: ""If you believe in science and that we have to act on climate change, then you have to vote!"" Hillary https://t.co/jfd"
nct_doyoungg|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
nct_doyoungg|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
_Dobbins_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
chicken_nuggit|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
chicken_nuggit|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
fcwic1|2ALAW|-0.5859|0.192|0.808|0.0|RT @2ALAW: Voter Fraud In PhiladelphiaPush Button One For HillaryPaid For By The Democratic County.#ElectionNight #DonaldTrump https:/
fcwic1||-0.5859|0.192|0.808|0.0|RT @2ALAW: Voter Fraud In PhiladelphiaPush Button One For HillaryPaid For By The Democratic County.#ElectionNight #DonaldTrump https:/
writingdownpat|ed_hooley|0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #ElectionDay #ElectionNight #Vote2016 #vote #USElection2016  https://t.
writingdownpat||0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #ElectionDay #ElectionNight #Vote2016 #vote #USElection2016  https://t.
darknessperrie|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
DrThomasPaul|DrThomasPaul|-0.8304|0.302|0.698|0.0|"RT @DrThomasPaul: #Hillary's extremely ill, evil and the most corrupt #politician the world may ever know. She's NOT for #America.#gmohttp"
hwomack2525|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
BelindaSpeight2|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
alison8796|Variety|0.0|0.0|1.0|0.0|RT @Variety: George W. Bush didn't vote for Donald Trump or Hillary Clinton for president https://t.co/JaXKzBWOTY https://t.co/CspXjAF5AS
alison8796|variety|0.0|0.0|1.0|0.0|RT @Variety: George W. Bush didn't vote for Donald Trump or Hillary Clinton for president https://t.co/JaXKzBWOTY https://t.co/CspXjAF5AS
BillyBobfagface|SophiaHelwani|0.6696|0.0|0.781|0.219|RT @SophiaHelwani: Hillary's greatest hits #7. Obama does the okie doke songl!  @placeboing @joerogan @TimKennedyMMA @Cowboycerrone @mitche
_ForeignStacks|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Nyro_LoL|OmniDestiny|0.1027|0.114|0.759|0.128|"RT @OmniDestiny: If Hillary wins and you're trying to get laid, there will probably be a lot of depressed Trumple chicks at the bars tonigh"
korbyn00|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Thats_Dessy|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
UdvTANBgkh9NQth|LuciaTaylor3|-0.4981|0.152|0.848|0.0|RT @LuciaTaylor3: @Suthen_boy There on the West side of Fl.  I passed 3 polling places and saw NO Hillary signs! #draintheswamp
thenatealdridge|HillaryforOH|0.5983|0.103|0.665|0.232|"RT @HillaryforOH: Rose escaped Nazi Germany at 15 &amp; is a proud American! Despite a recent broken hip, she just proudly cast her ballot for"
MaryEBarnes|DRUDGE_REPORT|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
MaryEBarnes|businessinsider|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
TheGoodGuy2016|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
turbo_thot_|drizzyxcole|0.5719|0.0|0.802|0.198|"RT @drizzyxcole: If Hillary wins Florida, do not slander my state for at least a week. https://t.co/skrGjKAgNl"
turbo_thot_|twitter|0.5719|0.0|0.802|0.198|"RT @drizzyxcole: If Hillary wins Florida, do not slander my state for at least a week. https://t.co/skrGjKAgNl"
SAILORSOLEMN|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
papiwhitelion|papiwhitelion|0.5719|0.0|0.812|0.188|RT @papiwhitelion: Will Bill Clinton be the 'First Man' of the USA if Hillary wins this Election?
mrsunshine44|AssangeFreedom|0.2481|0.092|0.761|0.146|RT @AssangeFreedom: @Wikileaks docs proved #Hillary seriously endangered  American security with her private email server! #ImVotingBecause
djwoolverton|PoliticsPeach|0.0|0.0|1.0|0.0|RT @PoliticsPeach: So the Bush Family didn't vote 4 Hillary Clinton after all... #ElectionNight
nosenseari|twitter|0.0|0.0|1.0|0.0|Cmon Hillary  #ImWithHer https://t.co/13CqFGjObn
Chloe2229|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
CLEFAlRlES|drewtoothpaste|0.4215|0.0|0.865|0.135|RT @drewtoothpaste: ME: anyone but trumpGARY JOHNSON: I will outlaw schools.JILL STEIN: Crystals are the only technology we need.ME: ok
TheSteveHolland|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
TheSteveHolland||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
aspen1031|blvckpapii|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
aspen1031|twitter|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
c_hallll|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
_hussonn|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
Dr__Bang|greeneyes0084|0.4215|0.0|0.882|0.118|"RT @greeneyes0084: #ImVotingBecause Hillary Clinton is the most corrupt person to ever seek the Presidency of the United States, &amp; she shou"
alexandraa2016|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
alexandraa2016|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Misty__Bella|Snapitson|0.3612|0.0|0.894|0.106|RT @Snapitson: Looks like #FBI agent that shot his wife..himself..burned down his house sent a message to #COMEY that was received loud &amp; c
dale_bernadette|seanhannity|-0.4574|0.187|0.813|0.0|@seanhannity Pennsylvania voters complained of their vote 2 Trump wld switch to Hillary. Frauding again?!
Kinara2_|Daniel_Oblak|-0.128|0.077|0.923|0.0|"@Daniel_Oblak I don't see any, and only one of the candidates has been caught trying to rig the elections. (Hillary)"
vexedmuddler|BitchestheCat|0.0|0.0|1.0|0.0|"RT @BitchestheCat: Every time a state gets called for Hillary, I'm doing a line of catnip. #ElectionDay https://t.co/kuqCiIhtLb"
vexedmuddler|twitter|0.0|0.0|1.0|0.0|"RT @BitchestheCat: Every time a state gets called for Hillary, I'm doing a line of catnip. #ElectionDay https://t.co/kuqCiIhtLb"
sunshinette|Pamela_Moore13|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
sunshinette|twitter|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
tsnkra|thetrudz|0.0|0.0|1.0|0.0|"RT @thetrudz: History, Symbolism &amp; Representation: Examining The Meaning of Hillary Rodham Clinton's Rise https://t.co/9EPPKpGgKe https://t"
tsnkra|thetrudz|0.0|0.0|1.0|0.0|"RT @thetrudz: History, Symbolism &amp; Representation: Examining The Meaning of Hillary Rodham Clinton's Rise https://t.co/9EPPKpGgKe https://t"
MattLegit10|LifeAsRednecks|0.6124|0.0|0.773|0.227|RT @LifeAsRednecks: Votin for Hillary just because shes a woman is like drinkin antifreeze just because it looks like Gatorade.
jimflynn39|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
tadiadunton|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
tadiadunton|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
JanetOmido|twitter|0.6145|0.0|0.555|0.445|YES! I VOTED FOR HILLARY CLINTON! https://t.co/fMjJ0mKuWU
VicColasanto|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
VicColasanto|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
NickStegmann|RowdyAmericans|0.0516|0.0|0.833|0.167|RT @RowdyAmericans: Hillary explained in 2 sentences https://t.co/nq0CsQIqBW
NickStegmann|twitter|0.0516|0.0|0.833|0.167|RT @RowdyAmericans: Hillary explained in 2 sentences https://t.co/nq0CsQIqBW
dihelfrich|tinkrbel5|-0.5106|0.125|0.875|0.0|RT @tinkrbel5: @DonaldJTrumpJr @Frankhe1 Right now I am sick of the soros owned machines recording Trump votes as Hillary in PA FL CA NC &amp;
anaxtaxhiamal|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
anaxtaxhiamal|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
curraheave|annalevinsonxx|-0.7739|0.226|0.774|0.0|"RT @annalevinsonxx: Im TIRED of this ""crooked Hillary"" rhetoric do u know how many times Donald has broken the law let GO of ur misogynY ht"
kimsgyeom|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
cherylmcfog|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
cherylmcfog|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
itsJustBClark|twitter|-0.34|0.103|0.897|0.0|"all over Facebook and it pisses me off, she goes on to say she voted for Hillary in the comments #podestaemails35 https://t.co/VtOyq1B116"
KameCobeEB|philsadelphia|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
KameCobeEB|twitter|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
VanessaLuver_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
VanessaLuver_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Sayitaintdaun|twitter|0.0|0.0|1.0|0.0|Is Hillary and Trump running still? https://t.co/13E4XJNOvo
skywolfangel|DilaChuu|-0.2755|0.297|0.703|0.0|RT @DilaChuu: I just don't like Hillary
Range2016|Pamela_Moore13|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
Range2016|twitter|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
zanesholtz|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
MY_PrettyAss|mefeater|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
MY_PrettyAss|twitter|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
hapihome|charliekirk11|0.4019|0.072|0.792|0.136|"RT @charliekirk11: Young voter and undecided? Watch this video: ""Hillary is part of the DC elite that has bankrupted America &amp; got rich o"
jlmcd13|JeffTutorials|0.3612|0.0|0.8|0.2|RT @JeffTutorials: .@HillaryClinton Just like you deleted your emails Crooked Hillary?
Barnett_59|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
pirateirwin|AFP|0.0|0.0|1.0|0.0|"RT @AFP: A large Hillary for America sign is displayed at the Jacob K. Javits Center in New York, where Clinton's #ElectionNight event is h"
Cuffs_No_Hoes|TheHomieLos|0.0|0.0|1.0|0.0|"RT @TheHomieLos: ""Vote for Hillary to keep Trump out of office""...I get it. But I need way more than that homie."
felicialindlov|itsellensalmon|0.0|0.0|1.0|0.0|RT @itsellensalmon: I know Hillary can do this! #ElectionNight
developertest09|twitter|0.0|0.0|1.0|0.0|Ouch for Hillary. Even if Indies only break for Trump +5% it would be OUCH. https://t.co/RqBOillxUd
UltralightBeth|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
UltralightBeth|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
_adornk|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_adornk|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
lgbtqtyIer|ridevocals|-0.4588|0.146|0.778|0.075|"RT @ridevocals: WHY ARE PEOPLE VOTING TRUMP BECAUSE ""HILLARY IS A CRIMINAL"" WHEN THE FBI ALREADY CLEARED HER AND TRUMP IS GOING TO COURT FO"
shyannesilvaa|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
shyannesilvaa|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
buckeyery|TattooedNnerdy|0.0|0.0|1.0|0.0|RT @TattooedNnerdy: #voted @TYTNetwork @HillaryClinton @realDonaldTrump #ElectionNight Hillary+Trump=  https://t.co/1BwijJ7flw
buckeyery|twitter|0.0|0.0|1.0|0.0|RT @TattooedNnerdy: #voted @TYTNetwork @HillaryClinton @realDonaldTrump #ElectionNight Hillary+Trump=  https://t.co/1BwijJ7flw
nellumbella|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
ymirius|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
ymirius|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
GuruVShetty|madhukishore|0.3612|0.0|0.848|0.152|RT @madhukishore: Like for Hillary or Retweet for Trump #ElectionDay #ElectionNight #ElectionFinalThoughts #USElection2016 #USADecides #Vot
__NaijaDrew|RUINER|-0.5719|0.381|0.619|0.0|"RT @RUINER: ""why do u hate Hillary?"" https://t.co/7fVEPi97U8"
__NaijaDrew|twitter|-0.5719|0.381|0.619|0.0|"RT @RUINER: ""why do u hate Hillary?"" https://t.co/7fVEPi97U8"
Tanner_hefner55|taebrooke|0.0|0.0|1.0|0.0|RT @taebrooke: All of Texas if Hillary is elected https://t.co/gPTQPVzZWx
Tanner_hefner55|twitter|0.0|0.0|1.0|0.0|RT @taebrooke: All of Texas if Hillary is elected https://t.co/gPTQPVzZWx
mikemyres12|AlGaldi|0.0|0.0|1.0|0.0|"RT @AlGaldi: #PresidentialElection sports comps.  I have #Trump as Steinbrenner, #Hillary as #ARod &amp; the race as a whole as the #MalaceAtTh"
acpcsn|voxdotcom|0.0|0.0|1.0|0.0|"Pantsuit Nation, the giant, secret Hillary Facebook group, explained https://t.co/MK06IlwK3A via @voxdotcom"
acpcsn|vox|0.0|0.0|1.0|0.0|"Pantsuit Nation, the giant, secret Hillary Facebook group, explained https://t.co/MK06IlwK3A via @voxdotcom"
jmay0418|twitter|0.0|0.0|1.0|0.0|This is the kind of woman Hillary thinks young women should listen to. #IvankaTrump is a class act compared to Mile https://t.co/wbB6Euke6j
alabaluu|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
alabaluu|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
BeccaRigal|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
PAClFRISK|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
PAClFRISK|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
goodforsumthin|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: Ohio, it's Election Day! Polls are open from 6:30am-7:30pm. Confirm your polling place now and go vote for Hillary! htt"
TheRogueelement|2ALAW|-0.4404|0.231|0.602|0.167|"RT @2ALAW: It's truly a sad day in America when we dismiss all the corruption, voting fraud committed as ""just politics""#Hillary is disqu"
DEE24_ALLStar|_Coca_cole_a|0.5719|0.0|0.748|0.252|RT @_Coca_cole_a: If Hillary wins I'll give everyone who rt's this $5
cutiepie9779|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
cutiepie9779|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
davidpwil|MissLizzyNJ|0.0|0.0|1.0|0.0|"RT @MissLizzyNJ: Remember, Hillary will take an early lead in exit polls which will change drastically, once Trump voters get out of work."
gnarruto|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
the_onlydime|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
LiamInfection|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
LiamInfection|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
MNVikingBeer|TheMorningSpew|0.3869|0.0|0.873|0.127|"RT @TheMorningSpew: Hillary is superstitious, so I thought we should cross her path with this: Please RT: @HillaryClinton #ElectionNight #M"
RipperBravoSix|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
fredgthegreat|halsteadg048|0.0|0.0|1.0|0.0|"RT @halsteadg048: Folks, in the two FL counties I've been watching, Hillary is DRAMATICALLY UNDERPERFORMING Obama.  We've got FL. https://t"
fredgthegreat||0.0|0.0|1.0|0.0|"RT @halsteadg048: Folks, in the two FL counties I've been watching, Hillary is DRAMATICALLY UNDERPERFORMING Obama.  We've got FL. https://t"
Gfabgab|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Gfabgab|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
annbeth22845|RichardGrenell|0.0|0.0|1.0|0.0|RT @RichardGrenell: Bridges in SoCal. Haven't seen anything for Hillary https://t.co/HCClZFt8eQ
annbeth22845|twitter|0.0|0.0|1.0|0.0|RT @RichardGrenell: Bridges in SoCal. Haven't seen anything for Hillary https://t.co/HCClZFt8eQ
BrookLassie|twitter|-0.7995|0.353|0.479|0.168|TOTALLY illegal.  hillary cheated in debate why wouldn't she steal an election? The woman had NO interest at her ra https://t.co/41jRUujXDG
JoshDavison024|FrankLuntz|0.6369|0.0|0.733|0.267|"RT @FrankLuntz: The numbers I'm getting now suggest a nationwide turnout that strongly favors Hillary.And if Hillary does well, so will d"
luvincowboys|DrThomasPaul|0.6114|0.0|0.81|0.19|RT @DrThomasPaul: Happy about this #LGBT/#LGBTQ for anyone who thinks #Hillary is for #gays? Think again!She's financing #murders.#gayhttp
peeltownembrys|twitter|-0.25|0.296|0.51|0.194|"Indeed, a Hillary win should scare the crap out of most foreigners. #warhawk https://t.co/lS52KXnmCa"
slendyisbae|Whathappen1d|0.3089|0.0|0.861|0.139|"RT @Whathappen1d: Americans, Harry very probably wants you to vote for Hillary, don't disappoint him"
s0phicee|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
s0phicee|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
jaira13s|FranchiseRocks|-0.9195|0.547|0.453|0.0|RT @FranchiseRocks: Damn bro. Hillary and Trump are the fucking devil. We're fucked.
Meguhhhh|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Meguhhhh|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
izzyfizzy1123|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
izzyfizzy1123|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
Paul55770744|linkis|0.9114|0.0|0.527|0.473|SEE IT! Madonna withdraws oral sex promise to Hillary voters https://t.co/nFe5tnhgGn. HA HA HA!! Have to watch video
pnam|twitter|-0.2755|0.117|0.883|0.0|Can't agree more Hillary will turn #US in to a corrupt banana republic Can't let that happen https://t.co/keXzYmsaFh
TheJMan91|SNFaizalKhamisa|0.327|0.0|0.872|0.128|@SNFaizalKhamisa why aren't we talking about the fact that Hillary deleted over a million emails??? ONE MILLION. Unbelievable.
hanxine|localblactivist|0.0|0.0|1.0|0.0|"RT @localblactivist: Similarly, Hillary has an infamous relationship with big money contributors."
brittytitty29|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
LeeLee_Ri|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
LeeLee_Ri|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
shanananananonn|brettt379|0.0772|0.0|0.86|0.14|RT @brettt379: I want 5 Valid reasons you voted for Hillary 
Lweendo23|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
heatherxstarrr|polaroidbones|-0.607|0.184|0.816|0.0|RT @polaroidbones: DONT SPLIT THE DEMOCRATIC VOTE TOMORROW CAUSE YOU DONT WANNA BE STUCK HILLARY OR TRUMP! ITS ONLY GONNA LEAVE US WITH TRU
Caam91|LiberalJaxx|-0.2263|0.173|0.722|0.105|RT @LiberalJaxx: I should have worn a hijab to vote for Hillary. Just to start some crap.  Getting my secret pleasures from the little thin
PlaidHeart|jkpresley|0.0|0.0|1.0|0.0|"RT @jkpresley: #ElectionNight *walks out of polling site*Reporter: ""how do you feel about just having voted for Hillary Clinton?""Me: htt"
moneeyy___|StahrMilan|-0.658|0.16|0.84|0.0|RT @StahrMilan: And to see people still down talking Hillary! Shut up bitch! When Bernie was running YALL ain't vote now it's Hillary and t
FCranmer|rorysutherland|-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
FCranmer||-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
Snikk|SLandinSoCal|0.0|0.0|1.0|0.0|RT @SLandinSoCal: Does #Hillary have #Kuru? Contracted through #Canabalism. Symptoms mimic #Parkinsons. Would explain her inappropriate out
ashley_hartage|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
SaBrown93|MicaBurton|0.4019|0.218|0.489|0.293|@MicaBurton i hope for your countries sake Hillary wins. no country should be burdened with Trump
throbbjon|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
blujaydavid|PerezHilton|0.0|0.0|1.0|0.0|RT @PerezHilton: #HillaryClinton does the #MannequinChallenge for #ElectionDay! https://t.co/EBHYc5eVrt https://t.co/i5Dz7zPnDo
blujaydavid|perezhilton|0.0|0.0|1.0|0.0|RT @PerezHilton: #HillaryClinton does the #MannequinChallenge for #ElectionDay! https://t.co/EBHYc5eVrt https://t.co/i5Dz7zPnDo
pedrobroa|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/GoYnDeEvaH
pedrobroa|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/GoYnDeEvaH
jazmineerae|___DestinyJadai|-0.6739|0.476|0.524|0.0|"RT @___DestinyJadai: ""VOTE HILLARY BITCH""  https://t.co/xVltWc6dU7"
jazmineerae|twitter|-0.6739|0.476|0.524|0.0|"RT @___DestinyJadai: ""VOTE HILLARY BITCH""  https://t.co/xVltWc6dU7"
yankeezag|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
marirodriguezim|lurrrveless|0.0|0.0|1.0|0.0|@lurrrveless Me too!! #imwithher #HillaryForPresident Go Hillary!! Go!! #GoVote
rhiannonbuquoii|WeekendSchemers|-0.3818|0.245|0.755|0.0|RT @WeekendSchemers: This is embarrassing. Hillary vs Hillary https://t.co/59K9hRKTe7
rhiannonbuquoii|twitter|-0.3818|0.245|0.755|0.0|RT @WeekendSchemers: This is embarrassing. Hillary vs Hillary https://t.co/59K9hRKTe7
carolineeileen_|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
carolineeileen_|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
S_Tiger_|sandkatt|-0.0276|0.227|0.552|0.221|RT @sandkatt: Can we really trust Hillary with the Chaos Emeralds?
nwonoway|TallahForTrump|0.1531|0.0|0.849|0.151|RT @TallahForTrump: How Hillary greets her corrupt little minions: https://t.co/4wn6HCASm6
nwonoway|twitter|0.1531|0.0|0.849|0.151|RT @TallahForTrump: How Hillary greets her corrupt little minions: https://t.co/4wn6HCASm6
Mr3lsewhere|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
Mr3lsewhere|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
jnblazz972|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
jnblazz972|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
deejjaaj|piercespears|0.5719|0.0|0.829|0.171|RT @piercespears: Historians will look back at this video and say this is why Hillary won the election  https://t.co/aaAKHIKPyv
deejjaaj|twitter|0.5719|0.0|0.829|0.171|RT @piercespears: Historians will look back at this video and say this is why Hillary won the election  https://t.co/aaAKHIKPyv
Push4Contest|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
jmw080|Autonomous138|0.3182|0.0|0.897|0.103|@Autonomous138 let us know how that 2% of the vote does in limiting the Democrat voter base Hillary's policies will expand.
BlastingNews|us|0.0|0.0|1.0|0.0|#election 2016 sees more #Facebook unfriending among #DonaldTrump and Hillary Clinton voters https://t.co/LfWSVgqUNR https://t.co/AfJAdNdbSU
kimlitwicki|TeamTrump|0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
kimlitwicki||0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
princejaygt|UglyGod|-0.5106|0.121|0.879|0.0|RT @UglyGod: It means yall shoulda fuckin listened &amp; kept Bernie Sanders as an option cause now we all look dumb af choosing between Hillar
Ebbi_Ling|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
valerie_orlando|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
indira_m9|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
constantino_sam|pinterest|-0.8208|0.457|0.543|0.0|TRUMP THAT BITCH - ANTI HILLARY PRO TRUMP POLITICAL BUMPER STICKER https://t.co/hlE23UztMY
mrobb1991|thenib|-0.049|0.113|0.784|0.103|"RT @thenib: ""I can't ignore that historically white feminism movements have ignored black and brown voices."" https://t.co/wHsFVaLS1A https:"
mrobb1991|thenib|-0.049|0.113|0.784|0.103|"RT @thenib: ""I can't ignore that historically white feminism movements have ignored black and brown voices."" https://t.co/wHsFVaLS1A https:"
iampicxsso|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
MattMolitov|WayneDupreeShow|-0.5754|0.189|0.811|0.0|RT @WayneDupreeShow: INSANE! PA Poll Workers Handing Out Instructions How To Vote For Hillary https://t.co/Pm1cBoHIoi #MyVote2016 #Election
MattMolitov|newsninja2012|-0.5754|0.189|0.811|0.0|RT @WayneDupreeShow: INSANE! PA Poll Workers Handing Out Instructions How To Vote For Hillary https://t.co/Pm1cBoHIoi #MyVote2016 #Election
GoddessOfTheOdd|Slate|0.5574|0.0|0.769|0.231|RT @Slate: Watch Hillary Clintons funniest off-script moments over 30 years: https://t.co/QrWHoKo5Je https://t.co/F22quZzObA
GoddessOfTheOdd|slate|0.5574|0.0|0.769|0.231|RT @Slate: Watch Hillary Clintons funniest off-script moments over 30 years: https://t.co/QrWHoKo5Je https://t.co/F22quZzObA
mallorykrenk|damnnnmoll|0.0|0.0|1.0|0.0|RT @damnnnmoll: I'd rather a cucumber be president instead of trump or hillary
DrThomasPaul|DrThomasPaul|0.4199|0.0|0.878|0.122|RT @DrThomasPaul: This #gay woman will tell you like it is. To the #gays brainwashed by #MSM: #WakeUP! #Hillary/#gmo #Trump #LGBTQhttps://
GeorgiaDaskalos|DRUDGE_REPORT|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
GeorgiaDaskalos|businessinsider|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
danarose1022|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
trapfentys|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
GetYouAStace|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
GetYouAStace|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
belly112|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
trenicole_|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
trenicole_|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Bethanygolatt|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Bethanygolatt|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
rstruglia17|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
rstruglia17|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
RealLifeChino|DonJuancho__|-0.2263|0.168|0.719|0.114|@DonJuancho__ true but no one wants Donald trump to become president. I'd rather Hillary
Kijwii|yvezayntIaurent|-0.5423|0.22|0.78|0.0|"RT @yvezayntIaurent: white person: idk whos worse: hillary or trumplgbtq, women, black people, immigrants, muslims: trump iswhite pers"
Smajor1995|AdamYT|0.9195|0.042|0.601|0.357|"@AdamYT @Seapeekay i find it so weird how like all the other states can vote trump, but if hillary gets like CA, NY, FL, WA, OH she wins ha"
GinoVelez201|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
kweenof_|twitter|0.0|0.0|1.0|0.0|#ivoted for Hillary Clinton #imwithher https://t.co/hEbYtPC5Vj
jammalama|FBI|0.0|0.0|1.0|0.0|"Conveniently, this news is too late. The @FBI should have been investing this weeks ago instead of reading more Hil https://t.co/hE9HpJOAUW"
jammalama|twitter|0.0|0.0|1.0|0.0|"Conveniently, this news is too late. The @FBI should have been investing this weeks ago instead of reading more Hil https://t.co/hE9HpJOAUW"
doobysnacks88|ShaySinches|0.0772|0.141|0.705|0.154|"@ShaySinches @brandiwilson318 hes not a politician and hes the perfect candidate, hillary though is a criminal and should not be running"
mhopson09|FortuneMagazine|0.7574|0.0|0.711|0.289|honoring those who came before you! Why Hillary Clinton supporters are wearing white to vote via @FortuneMagazine https://t.co/0LFUXAgnaW
mhopson09|fortune|0.7574|0.0|0.711|0.289|honoring those who came before you! Why Hillary Clinton supporters are wearing white to vote via @FortuneMagazine https://t.co/0LFUXAgnaW
theriseofgomez|vibeeeez|-0.5574|0.261|0.739|0.0|RT @vibeeeez: prediction: Hillary Clinton is our next present &amp; everyone is shocked Trump lost
choiteas|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
choiteas|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
Upsunson|DVATW|0.5106|0.0|0.87|0.13|RT @DVATW: Bill Clinton tried to cheer up Hillary today by reminding her that Mandela wasn't elected president until after serving 27 yrs i
youngbola1|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Gem_Crazy_81|BunaTime|-0.5859|0.174|0.826|0.0|"RT @BunaTime: ""When zat bitch Hillary takes over, you can come here anytime and drink buna with us"" https://t.co/KcvvS4s8sW"
Gem_Crazy_81|twitter|-0.5859|0.174|0.826|0.0|"RT @BunaTime: ""When zat bitch Hillary takes over, you can come here anytime and drink buna with us"" https://t.co/KcvvS4s8sW"
angellbadass|BalmainBoslick|-0.1027|0.065|0.935|0.0|RT @BalmainBoslick: Everybody keep askin who I'm voting for idk Hillary gon take my Guns &amp; Trump gon take my FoodStamps
rharrisonfries|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana 0.5% reporting TRUMP 70.1% | Hillary 26.1% massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Electi
ItzKurisu|bawbbyspears|0.5106|0.0|0.852|0.148|RT @bawbbyspears: Fun fact: Britney Spears was Hillary's first choice for Vice President. Britney declined because she's a mom now. https:/
ItzKurisu||0.5106|0.0|0.852|0.148|RT @bawbbyspears: Fun fact: Britney Spears was Hillary's first choice for Vice President. Britney declined because she's a mom now. https:/
Angelmdunn1961|zachhaller|0.5267|0.0|0.784|0.216|RT @zachhaller: Hillary is a straight up robot.She legit needs handlers to remind her to act like a human.#PodestaEmails33/52567 https:
brockheather03|JackPosobiec|-0.2023|0.141|0.859|0.0|RT @JackPosobiec: LIVE on #Periscope: Hillary Workers Intimidate Voters in Philly https://t.co/u9aM89xnPY
brockheather03|periscope|-0.2023|0.141|0.859|0.0|RT @JackPosobiec: LIVE on #Periscope: Hillary Workers Intimidate Voters in Philly https://t.co/u9aM89xnPY
Aprado7997|riyasharma266|0.1779|0.14|0.667|0.194|RT @riyasharma266: Remember those four brave men who asked Hillary for help 700 times before they were murdered. Think of them on VOTING DA
Dre_NoOvO|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
wavvycee|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
wavvycee|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
rachel_obrien14|PriceAbby1|0.0|0.0|1.0|0.0|"RT @PriceAbby1: I think the first 33,000 votes for Hillary should get deleted right?"
Didnttii|TheWorldOfFunny|0.0|0.0|1.0|0.0|RT @TheWorldOfFunny: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/rYVq0sC4U5
Didnttii|twitter|0.0|0.0|1.0|0.0|RT @TheWorldOfFunny: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/rYVq0sC4U5
Harley_Woody|uproxx|0.0258|0.112|0.769|0.118|"If Youre Still Undecided, Let These Rappers Convince You To Vote For Hillary Clinton https://t.co/lzPrnxMCH1"
braxtonmasters_|Sadieisonfire|0.2732|0.138|0.667|0.195|RT @Sadieisonfire: damn I can't believe this was the deciding factor that made Hillary win https://t.co/tEo4vvVmNj
braxtonmasters_|twitter|0.2732|0.138|0.667|0.195|RT @Sadieisonfire: damn I can't believe this was the deciding factor that made Hillary win https://t.co/tEo4vvVmNj
sarahimages|nytimes|0.0|0.0|1.0|0.0|Life in the Lights https://t.co/QODdFFqpJ0
NoBrakesAndrew|Jawwwwwsh|0.5719|0.0|0.817|0.183|RT @Jawwwwwsh: Vote for Hillary so we can experience the Tomi Lahren mental breakdown. That entertainment is worth more than the future of
lildolcezza|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
tamaraleighllc|KingAJ40|0.6209|0.0|0.747|0.253|RT @KingAJ40: Good People of UTAH!!! Don't Let Hillary Clinton CONFISCATE your GUNS!!!https://t.co/E7zbgg966nhttps://t.co/I97WEXYJNE
tamaraleighllc|t|0.6209|0.0|0.747|0.253|RT @KingAJ40: Good People of UTAH!!! Don't Let Hillary Clinton CONFISCATE your GUNS!!!https://t.co/E7zbgg966nhttps://t.co/I97WEXYJNE
Giannaamarieeee|owensupertramp|0.2105|0.256|0.407|0.338|RT @owensupertramp: don't mistake my hate for trump with support for hillary. we're either fucked or super weenie hut fucked
wworkergates|GovMikeHuckabee|0.0|0.0|1.0|0.0|"RT @GovMikeHuckabee: State Dept says it takes 5 yrs to review 31,000 Hillary emails. Let Comey do it!  He can review 650,000 in 1 week!  ht"
vyntage_lo|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
vyntage_lo|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
mahabouraoud|Team_Smoldy|0.0|0.0|1.0|0.0|@Team_Smoldy @CherylH64579178 @iansomerhalder an hour later Hillary would call him and say come to the office. She made a lot of Bill's
CLEFAlRlES|drewtoothpaste|0.0|0.0|1.0|0.0|"RT @drewtoothpaste: And in our final debate, the third pa-BILL WELD: Vote for Hillary.GARY JOHNSON: He didn't say that. Fake.JILL STEIN:"
Sesh_Jayy|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Sesh_Jayy|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
haleyhauskins|ShouldersTaylor|0.34|0.0|0.861|0.139|RT @ShouldersTaylor: I want to get married. And have kids. And live my life. And I believe if Hillary becomes president God will end this w
michaelvlueder|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
michaelvlueder|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
kihyanaee|Amxlorde|0.7269|0.0|0.736|0.264|RT @Amxlorde: look I just pray that Hillary win tonight  if not we gone need to come together as a whole 
Courtney_Mackk|TheOneandOnIyUS|0.7096|0.0|0.753|0.247|RT @TheOneandOnIyUS: The joke is on Hillary if she wins. She'll have to sit at the desk Monica sat under.
RealJoeMirto|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
VEN0MKlNG|GraphicTweetss|-0.6124|0.364|0.636|0.0|RT @GraphicTweetss: Trump = open racistHillary = closet racist https://t.co/6QK3XJe2ID
VEN0MKlNG|twitter|-0.6124|0.364|0.636|0.0|RT @GraphicTweetss: Trump = open racistHillary = closet racist https://t.co/6QK3XJe2ID
Sammmyyy_25|brookeregalado|0.8276|0.0|0.734|0.266|"RT @brookeregalado: if you vote for hillary &amp; she wins, you better not complain when the U.S. goes down in flames bc you're the one that ga"
Virtualnsainity|ltsDonaIdTrump_|0.0|0.0|1.0|0.0|RT @ltsDonaIdTrump_: Hillary Clinton's da sells avon
RealJobRob|bad_bad_bernie|-0.1828|0.148|0.738|0.114|RT @bad_bad_bernie: It wasn't the Republicans attacking Hillary that destroyed the Democratic Party.It was the Democrats defending Hillar
Natalienikole_|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Natalienikole_|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
kategoellerr|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
kategoellerr|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
braedontalley|JLaughmiller|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
braedontalley|twitter|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
Kent_Cyclist|D_Blanchflower|0.0|0.0|1.0|0.0|RT @D_Blanchflower: The name Trump should from this day forward be synonymous with everything we teach our children not to become... 1/2ht
ElHombreBDD|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
DLPaxt|AtlTeaPartyLove|0.0|0.0|1.0|0.0|"RT @AtlTeaPartyLove: If your Role Models are Jay Z, Beyonce and GaGa. You voted for Hillary because they told you to. Then, you already los"
SelfMade_Tye|GIRLHEFUNNY|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
SelfMade_Tye|twitter|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
monicapaos|Laughbook|0.0|0.0|1.0|0.0|RT @Laughbook: When you have to vote for Trump or Hillary #ElectionDay https://t.co/NKBZfMN4Ys
monicapaos|twitter|0.0|0.0|1.0|0.0|RT @Laughbook: When you have to vote for Trump or Hillary #ElectionDay https://t.co/NKBZfMN4Ys
vincesaiz1|theScore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
vincesaiz1|thescore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
spnsammy|patrickhumps|-0.4588|0.19|0.724|0.086|RT @patrickhumps: If Hillary loses the election by like 1 vote I'm blaming it on the person who wrote in Harry Styles on their ballot
Eric_Dockery1|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Polysexuals|tugbeck|0.0268|0.3|0.433|0.267|"RT @tugbeck: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost. #ElectionDay"
Williamrmontgo1|DonaldJTrumpJr|-0.3229|0.179|0.737|0.084|@DonaldJTrumpJr that is very true Hillary will not protect this country she might sell it out but she won't protect it
geena1017|mefeater|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
geena1017|twitter|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
OfficalHillary|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
DorH84607784|LeighPatrick|0.0|0.0|1.0|0.0|"RT @LeighPatrick: Given the reports flooding in nationwide, you either vote Hillary or the machine votes Hillary for you. #Corruption #elec"
SaraiCruz10_|ClarenceJWhite|0.0|0.069|0.863|0.069|RT @ClarenceJWhite: I feel like Trump &amp; Hillary are two divorced parents fighting over custody of us but we kinda just wanna go live with g
gpreudhomme|DavidCornDC|0.0|0.0|1.0|0.0|RT @DavidCornDC: Where Hillary Clinton will declare victory or....something else. https://t.co/4b82Lt4UGB
gpreudhomme|twitter|0.0|0.0|1.0|0.0|RT @DavidCornDC: Where Hillary Clinton will declare victory or....something else. https://t.co/4b82Lt4UGB
leinani_cambra|stein_baraka|0.0|0.0|1.0|0.0|RT @stein_baraka: #ElectionDay #PopQuiz: Hillary Clinton is....#jillnothill #podestaemails35 #maga #imwithher #ivoted #poll #jillstein201
donna_grooms|TIME|-0.0258|0.073|0.927|0.0|RT @TIME: The overlooked history behind the movement to wear white on Election Day https://t.co/4aYW2SdOcG
donna_grooms|time|-0.0258|0.073|0.927|0.0|RT @TIME: The overlooked history behind the movement to wear white on Election Day https://t.co/4aYW2SdOcG
Ziii_10|Chico_Mills|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
Ziii_10|twitter|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
FallingAngel790|DESlRABLE|-0.533|0.194|0.723|0.084|@DESlRABLE @Calum5SOS definitely not Jesus 2.0 but I'm more scared of what Hillary will do compared to Trump
Shelby_999_|porn_horse|-0.7656|0.292|0.708|0.0|RT @porn_horse: Hillary campaigner employed FORBIDDEN MAGIC to do a kickflip in heels. No one is talking about this!!!https://t.co/GD9L0u
Shelby_999_|t|-0.7656|0.292|0.708|0.0|RT @porn_horse: Hillary campaigner employed FORBIDDEN MAGIC to do a kickflip in heels. No one is talking about this!!!https://t.co/GD9L0u
Annie_lovessPR|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
lmkwhitesides|ridevocals|-0.4588|0.146|0.778|0.075|"RT @ridevocals: WHY ARE PEOPLE VOTING TRUMP BECAUSE ""HILLARY IS A CRIMINAL"" WHEN THE FBI ALREADY CLEARED HER AND TRUMP IS GOING TO COURT FO"
NickBent|rorysutherland|-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
NickBent||-0.5994|0.151|0.849|0.0|RT @rorysutherland: Fact: Hillary Clinton would be the first female American head of state since the death of Queen Anne in 1714. https://t
alexschickel|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
babyyogy1964|BillHemmer|0.4576|0.0|0.75|0.25|@BillHemmer @HillaryClinton @realDonaldTrump I think Trump is more trusting then hillary
Sq0410|OhNoSheTwitnt|0.4168|0.0|0.883|0.117|RT @OhNoSheTwitnt: Out to dinner in North Carolina wearing my Hillary shirt. It's under a sweater though I'm not stupid these people have g
sharpinkner|pizzaparacenar|0.0|0.0|1.0|0.0|RT @pizzaparacenar: Ni Trump ni Hillary https://t.co/O4X2zybhAX
sharpinkner|twitter|0.0|0.0|1.0|0.0|RT @pizzaparacenar: Ni Trump ni Hillary https://t.co/O4X2zybhAX
SlinkysAfreak|Slate|0.5574|0.0|0.769|0.231|RT @Slate: Watch Hillary Clintons funniest off-script moments over 30 years: https://t.co/QrWHoKo5Je https://t.co/F22quZzObA
SlinkysAfreak|slate|0.5574|0.0|0.769|0.231|RT @Slate: Watch Hillary Clintons funniest off-script moments over 30 years: https://t.co/QrWHoKo5Je https://t.co/F22quZzObA
tlvrp_russia|therussophile|-0.6597|0.206|0.794|0.0|#Moscow #SaintPetersburg Proof That 100 Years of Voting for the Lesser Evil Gave Us Trump and Hillary https://t.co/Vzqd2EPmbp
JR777771|kindcutesteve|-0.5719|0.209|0.791|0.0|RT @kindcutesteve: MotherJones: This Election Is a Referendum on Hate (vote against it)#p2 #TNTweeters #USLatino #VoteBluehttps://t.co/Yj
TheMource|themource|0.2755|0.0|0.869|0.131|for more info https://t.co/6fXFivzEre Hillary Clinton -- Don't Mess W... https://t.co/nEp8eeyHqw #lol #cute #live https://t.co/EBi78lXDYa
_gloooooria|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_gloooooria|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
dotsmack|LisaClaire9090|0.3973|0.0|0.871|0.129|"RT @LisaClaire9090: @Anne_Nissell @dotsmack We MUST Include Our #WestCoast Americans, as Far West as #Hawaii Final Count Very Important!! W"
Charlamaigne|HaskelBiz|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
Charlamaigne|twitter|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
Danieljackson94|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
Danieljackson94|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
eurekajimbob|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
JimSjim409|Cubs|0.6597|0.109|0.565|0.327|"God, Said I wouldnt ask for anything for awhile since the @Cubs won but.....Lord, Please let Hillary lose. OH...AMEN"
Nighthawkrlder|OnlineMagazin|-0.5267|0.207|0.714|0.079|RT @OnlineMagazin:  That made my day. Crooked Hillary supporter went into the trap when he wanted to steal the #DonaldTrump shield. ht
ikeaah|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
_kayaleigh_|MorganSchuette|-0.6166|0.366|0.634|0.0|RT @MorganSchuette: TRUMP FOR PRESIDENT HILLARY FOR PRISON
wingate_david|CNN|0.0|0.0|1.0|0.0|@CNN @HillaryClinton @realDonaldTrump We all know the journalists at #CNN are on HILLARY'S payroll.I will pass on watching you.#TrumpTV
FreeUs551|DrThomasPaul|0.3612|0.0|0.878|0.122|"RT @DrThomasPaul: This sums you up #Obama. 97 to 1 agree. Obama/#Hillary, You're not #Americans. #Trump #Bernie #Sept11 #Election2016 https"
KelsoOConnor|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
Creekredman|worldnetdaily|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
Creekredman|wnd|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
Deserie_Larios|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Deserie_Larios|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
SincerelyWendy|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
ctimm75|emmavanalstine9|0.0|0.0|1.0|0.0|RT @emmavanalstine9: Anyone but Hillary
Alexiaa_Minaj|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
ladykatrina3|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
ladykatrina3|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
_BigBobbyD_|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
_BigBobbyD_|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
i_wokeuplikedis|bigshitxtalker|0.0|0.0|1.0|0.0|RT @bigshitxtalker: Polls close at 7 pm. Hurry up and get in line and vote for Hillary. https://t.co/rBZu2LjQlJ
i_wokeuplikedis|twitter|0.0|0.0|1.0|0.0|RT @bigshitxtalker: Polls close at 7 pm. Hurry up and get in line and vote for Hillary. https://t.co/rBZu2LjQlJ
s5xfast|WhitePeepsDo|-0.4767|0.255|0.745|0.0|"RT @WhitePeepsDo: Forget Trump and Hillary, this man Gary Johnson has no chill https://t.co/c5nOgggTd8"
s5xfast|twitter|-0.4767|0.255|0.745|0.0|"RT @WhitePeepsDo: Forget Trump and Hillary, this man Gary Johnson has no chill https://t.co/c5nOgggTd8"
CallOfBeautyy_|GIRLHEFUNNY|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
CallOfBeautyy_|twitter|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
tljbd|Scarlett210|-0.765|0.28|0.72|0.0|"RT @Scarlett210: And #Hillary is a self-serving #elitist who'll continue #globalist policies, destroy ur safety&amp; deprive ur kids of a futur"
Casmir_Egbe|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
Casmir_Egbe|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
61Rinaldi|JoshuaThifault|-0.38|0.237|0.626|0.137|RT @JoshuaThifault: Hillary trying to steal Florida!! Is anyone really surprised? https://t.co/dGahBpE8VH
61Rinaldi|twitter|-0.38|0.237|0.626|0.137|RT @JoshuaThifault: Hillary trying to steal Florida!! Is anyone really surprised? https://t.co/dGahBpE8VH
Smedley_Butler|ActualFlatticus|-0.6908|0.207|0.793|0.0|"RT @ActualFlatticus: We already do that.  Obama, and specifically Panetta, who Hillary will be appointing to something, intentionally kill"
memotaur|ReturnofRV|0.1779|0.109|0.746|0.144|"RT @ReturnofRV: Why are all the Hillary supporters, Hillary trolls, and Hillary mainstream media pundits strangely quiet?"
teri3626|BreitbartNews|0.2924|0.299|0.289|0.413|@BreitbartNews Hillary wonderful voters! Gross!
todd_anuchitN|theScore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
todd_anuchitN|thescore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
peachymarz|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
JayC2x|GIRLHEFUNNY|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
JayC2x|twitter|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
AllLivesMtr81|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
tweetwithtee|marwannafuq|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
tweetwithtee|twitter|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
SaskiaHallenga|FrankLuntz|0.6369|0.0|0.733|0.267|"RT @FrankLuntz: The numbers I'm getting now suggest a nationwide turnout that strongly favors Hillary.And if Hillary does well, so will d"
twosontribune|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
twosontribune|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
tee_shelton|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
tee_shelton|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
a_cosgrove|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
kelly_heroes|PrinceRoyce|0.5719|0.0|0.619|0.381|@PrinceRoyce Hillary loves his little man bun
BrittanyFlore16|TheChainsmokers|0.0|0.0|1.0|0.0|RT @TheChainsmokers: lets get a little early chainsmoker election poll going... Trump or Hillary... vote below
InOtherNewsNotO|AssangeFreedom|0.4559|0.058|0.797|0.145|RT @AssangeFreedom: #ImVotingBecause Its my duty to clean corruption out of my country! @Wikileaks exposed #Hillary with her OWN documents!
Nola_Darling84|ShaanMKhan|0.0|0.0|1.0|0.0|RT @ShaanMKhan: Hillary Clinton's platform includes $25 Billion for HBCUs! Let's ELECT HER and hold her ACCOUNTABLE! Don't forget!#Electi
chickensherri|ThatSusanBurke|-0.1531|0.071|0.929|0.0|RT @ThatSusanBurke: Tomorrow Hillary will start planning her presidency and Trump will file lawsuits &amp; figure out products for his new luxu
DamnGirlMelanie|mefeater|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
DamnGirlMelanie|twitter|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
pfunbun|ptownjake|0.3804|0.0|0.844|0.156|RT @ptownjake: Very cool. #Portland music licensing company @marmosetmusic curated Hillary's campaign playlist. #imwithher https://t.co/C9b
pfunbun|t|0.3804|0.0|0.844|0.156|RT @ptownjake: Very cool. #Portland music licensing company @marmosetmusic curated Hillary's campaign playlist. #imwithher https://t.co/C9b
_sogofiez|officialSmith_|0.3612|0.0|0.783|0.217|RT @officialSmith_: *casts vote for Hillary*Hillary: Thank you s--Me: https://t.co/rmDqKBTo1i
_sogofiez|twitter|0.3612|0.0|0.783|0.217|RT @officialSmith_: *casts vote for Hillary*Hillary: Thank you s--Me: https://t.co/rmDqKBTo1i
brady_benner|officialSmith_|0.3612|0.0|0.783|0.217|RT @officialSmith_: *casts vote for Hillary*Hillary: Thank you s--Me: https://t.co/rmDqKBTo1i
brady_benner|twitter|0.3612|0.0|0.783|0.217|RT @officialSmith_: *casts vote for Hillary*Hillary: Thank you s--Me: https://t.co/rmDqKBTo1i
junecrotty|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
jaydaSlays|PETTYMAMII|-0.8441|0.269|0.731|0.0|RT @PETTYMAMII: Vote Hillary Clinton idc is she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
freeandfunny14|NewsweekEurope|0.0|0.0|1.0|0.0|RT @NewsweekEurope: Read Julian Assange's statement on why Wikileaks has published Clinton campaign documents https://t.co/ojoq2RmEpV https
freeandfunny14|newsweek|0.0|0.0|1.0|0.0|RT @NewsweekEurope: Read Julian Assange's statement on why Wikileaks has published Clinton campaign documents https://t.co/ojoq2RmEpV https
EsKearl|theScore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
EsKearl|thescore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
Lord_Sebastian3|Cali_Kid_7|-0.296|0.167|0.833|0.0|RT @Cali_Kid_7: If Hillary gets elected I'm moving to Benghazi... at least I know she'll leave me alone there..
stonadarico|marwannafuq|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
stonadarico|twitter|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
erreavecmoi|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
erreavecmoi|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
gatitadelrey|arzE|0.7865|0.0|0.729|0.271|RT @arzE: voting for Hillary doesn't have to be ur longest yeah boy ever. It can be ur shorter yeah boy ever. Just uhh don't waste ur yeah
catalinanemmi|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
suhasinih|AFP|0.0|0.0|1.0|0.0|"RT @AFP: A large Hillary for America sign is displayed at the Jacob K. Javits Center in New York, where Clinton's #ElectionNight event is h"
mariajoao2101|Chico_Mills|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
mariajoao2101|twitter|0.3612|0.0|0.737|0.263|RT @Chico_Mills: Like For TrumpRetweet For Hillary https://t.co/Ab6MfMWlAd
Logan41114743|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Logan41114743|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Amituofo2013|NewsPho|0.0|0.0|1.0|0.0|RT @NewsPho: @Breaking911 Voting Machines #Rigged for Hillary Clinton. #VoterFraud #ElectionDay #USelection2016 https://t.co/6lkJ9n1U8R
Amituofo2013|twitter|0.0|0.0|1.0|0.0|RT @NewsPho: @Breaking911 Voting Machines #Rigged for Hillary Clinton. #VoterFraud #ElectionDay #USelection2016 https://t.co/6lkJ9n1U8R
Luckyyou__|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Luckyyou__|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
RedotZone|redotzone|0.4019|0.0|0.769|0.231|Rihanna Wears Her Support for Hillary Clinton Again https://t.co/3p1goZYxzB https://t.co/ybz9FyWqzw
megannn_23|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
carmonyj34|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
carmonyj34|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
cam6499|cristinalaila1|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
cam6499|twitter|0.0|0.0|1.0|0.0|"RT @cristinalaila1: Trump has 251,000 Retweets vs Hillary's 32,000 and she even pinned  her tweet #ElectionDay https://t.co/EV1LJPn1wg"
Bennzie|KatiCut|-0.8142|0.271|0.729|0.0|@KatiCut Hillary is a vote for more of the same corrupt bullshit. Trump is a vote for change. Absolutely not the 2 greatest candidates tho..
CallistroFlores|Things4Guys|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
CallistroFlores|twitter|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
judediab2|Oldfirmfacts1|0.0|0.0|1.0|0.0|"RT @Oldfirmfacts1: Trump: ""Hillary must release the 33,000 emails""Celtic matchday announcer: ""Yeah, release the 56,412 emails"""
_nne_nne|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
NikoMarcella|JohnnyWojo|0.743|0.0|0.76|0.24|"RT @JohnnyWojo: If Hillary wins, I'm moving to Mexico and then sneaking back into the US so I can reap all the benefits."
JSara1234|mikethenice1|0.1779|0.0|0.866|0.134|RT @mikethenice1: BREAKING: Latest National Polls Show Trump With Growing Lead https://t.co/H3SoiijcM9
JSara1234|conservativetribune|0.1779|0.0|0.866|0.134|RT @mikethenice1: BREAKING: Latest National Polls Show Trump With Growing Lead https://t.co/H3SoiijcM9
roxy6118|worldnetdaily|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
roxy6118|wnd|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
Kykylaaaaaa|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Kykylaaaaaa|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
UdvTANBgkh9NQth|Suthen_boy|0.0|0.0|1.0|0.0|RT @Suthen_boy: This is at a polling station in Ft Lauderdale FL - not a single Hillary sign.    #tcot #ccot #MAGA #draintheswamp https://t
UdvTANBgkh9NQth||0.0|0.0|1.0|0.0|RT @Suthen_boy: This is at a polling station in Ft Lauderdale FL - not a single Hillary sign.    #tcot #ccot #MAGA #draintheswamp https://t
kailacamillia|jesieraybrown|-0.521|0.325|0.675|0.0|RT @jesieraybrown: #ImVotingBecause  we can't let Hillary win!
TheBigToenail|Mike3453Mike|-0.4588|0.131|0.805|0.064|RT @Mike3453Mike: Is this why Marines die. That is to say to allow Hillary Clinton's rise as did Hitler to be above a Nation's rule of law.
5SOSWWReports|melina312_|0.5719|0.0|0.575|0.425|@melina312_ Even if Hillary wins tho
eli_arza|dfernandezz_|-0.92|0.389|0.611|0.0|RT @dfernandezz_: Bitch said she can't vote for Hillary cause she's a liar YOUR MAN'S A LIAR AND YOU'RE STILL WITH HIM SO ???????
Idolme922|MrDane1982|0.0|0.0|1.0|0.0|RT @MrDane1982: Little kids walking through Harlem chanting vote!!!! I'm with Hillary Clinton! https://t.co/haAlItIYzT
Idolme922|twitter|0.0|0.0|1.0|0.0|RT @MrDane1982: Little kids walking through Harlem chanting vote!!!! I'm with Hillary Clinton! https://t.co/haAlItIYzT
clifjules|money|0.0|0.0|1.0|0.0|"George W. Bush did not vote for Clinton, despite what Rush Limbaugh claimed https://t.co/iJFHvH3BwT #online"
DanielRicciulli|FiveThirtyEight|0.5859|0.0|0.798|0.202|"According to @FiveThirtyEight prediction, Hillary Clinton is set to win with a 71% majority over Donald Trump"
Buffy619|extratv|0.3818|0.0|0.809|0.191|RT @extratv: Would @CoryBooker accept a position in a @HillaryClinton cabinet? https://t.co/SaGHTasbXe #ElectionDay https://t.co/xV8a2h6RqF
Buffy619|extratv|0.3818|0.0|0.809|0.191|RT @extratv: Would @CoryBooker accept a position in a @HillaryClinton cabinet? https://t.co/SaGHTasbXe #ElectionDay https://t.co/xV8a2h6RqF
janismclaren1|mitchellvii|0.4404|0.0|0.861|0.139|RT @mitchellvii: I'm noticing the exit polls from MSNBC are dramatically better for Hillary than the ones from Fox.
KeepItTricky|LouisFarrakhan|0.7579|0.0|0.683|0.317|@LouisFarrakhan @joeyBADASS glad to see someone hasn't sold their soul to Hillary's false sense of optimism.
_fossit_|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
_fossit_|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
KDay1937|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
richsp8jr|LosEddy|0.1901|0.0|0.907|0.093|"RT @LosEddy: Mexicans today are all like ""Go Hillary you got this"" but on Friday.. ""VIVA MEXICO CABRONES"" "
sonjamart48|US_Army_Vet|0.0|0.0|1.0|0.0|RT @US_Army_Vet: Hillary had her maid print classified mat'l: NYPhttps://t.co/lEur7MncMo Breitbarthttps://t.co/q2nerd6kVU @American1765 @
icyforoccasion|pieceofjay|0.0|0.0|1.0|0.0|RT @pieceofjay: JUST FUCKING VOTE FOR HILLARY
nellyaandalon|GIRLHEFUNNY|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
nellyaandalon|twitter|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
seanwlknsn|Americooligan|0.0|0.0|1.0|0.0|"RT @Americooligan: Trump up 70.5% to Hillary's 25.8% in Indiana. 35,646 votes to 13,049 (1% reporting). #ElectionNight"
IdkGoAskYourMom|HoltBlack05|-0.4404|0.367|0.633|0.0|RT @HoltBlack05: Hillary Clinton hates puppies
APikeGoff|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
APikeGoff|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
_Smilerzxx|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
_Smilerzxx|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Lnkobin|twitter|-0.5423|0.226|0.774|0.0|Fuck Hillary&amp;Trump my nigga Stone Cold got my vote all the waaay  https://t.co/XuMZROylhd
ReligionRetards|TaShanna10|0.6908|0.0|0.778|0.222|@TaShanna10 Hillary is using U for a vote again &amp; will not bring jobs or opportunity. She is good at laundering money to ClintonFoundation.
texasmfg|weknowwhatsbest|-0.2263|0.139|0.759|0.101|RT @weknowwhatsbest: President Obama endorses Hillary because she's the only candidate who has experience in carrying out his failed polici
Tigers930410|jaynordlinger|0.7579|0.0|0.745|0.255|"RT @jaynordlinger: Hillary = luckiest politician ever. I know the hour is late, but are we SURE that Trump was not a Clinton plant?"
kysgabbygirl|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
Korizwick|DontTread_2nd|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
Korizwick|twitter|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
amatangy|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
jbyrons83|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
_Jaedore|ASAP_Toby|0.296|0.0|0.784|0.216|@ASAP_Toby a joke for a woman to become president or Hillary ?
VedehiMajumdar|kylegriffin1|0.5267|0.0|0.804|0.196|RT @kylegriffin1: Inbox: Hillary for America Statement in Support of Bipartisan Efforts to Extend Voting Hours in Durham County. https://t.
VedehiMajumdar||0.5267|0.0|0.804|0.196|RT @kylegriffin1: Inbox: Hillary for America Statement in Support of Bipartisan Efforts to Extend Voting Hours in Durham County. https://t.
torijudah|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
torijudah|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
DragemT1814|marwannafuq|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
DragemT1814|twitter|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
tayelurade|sadgallexi|-0.5106|0.142|0.858|0.0|"RT @sadgallexi: ""Hillary is a liar, listen to me while I parrot things people have been saying for years to sound smart."" https://t.co/sN2A"
tayelurade|t|-0.5106|0.142|0.858|0.0|"RT @sadgallexi: ""Hillary is a liar, listen to me while I parrot things people have been saying for years to sound smart."" https://t.co/sN2A"
Hunter_Ash23|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
gracelongg_|mykebm|-0.09|0.119|0.779|0.101|"RT @mykebm: idc Hillary is better than trump , I mean they're both shit but u gotta weigh your options"
drdonna212|CNN|-0.3382|0.23|0.77|0.0|@CNN I think Comey voted for Hillary out of guilt!
judithshaw2|worldnetdaily|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
judithshaw2|wnd|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
lolkiyaa|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
lolkiyaa|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
Jatyrz|huffpostqueer|0.4404|0.0|0.818|0.182|RT @huffpostqueer: Here's why Hillary Clinton supporters stormed the Brooklyn Bridge in pantsuits https://t.co/3vM07ezKXp
Jatyrz|huffingtonpost|0.4404|0.0|0.818|0.182|RT @huffpostqueer: Here's why Hillary Clinton supporters stormed the Brooklyn Bridge in pantsuits https://t.co/3vM07ezKXp
WhiskeyStr8Up|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
WhiskeyStr8Up|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
G_isellegomez|LosEddy|0.1901|0.0|0.907|0.093|"RT @LosEddy: Mexicans today are all like ""Go Hillary you got this"" but on Friday.. ""VIVA MEXICO CABRONES"" "
_enrolandote|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
larus_minutus|ActualFlatticus|-0.765|0.248|0.752|0.0|RT @ActualFlatticus: Has Hillary Clinton ever said a single word that led you to believe she intends to stop killing people in 7 countries?
peepmyprogress|Slate|0.5574|0.0|0.769|0.231|RT @Slate: Watch Hillary Clintons funniest off-script moments over 30 years: https://t.co/QrWHoKo5Je https://t.co/F22quZzObA
peepmyprogress|slate|0.5574|0.0|0.769|0.231|RT @Slate: Watch Hillary Clintons funniest off-script moments over 30 years: https://t.co/QrWHoKo5Je https://t.co/F22quZzObA
Toni18000954|navyseal6|-0.6808|0.189|0.811|0.0|"RT @navyseal6: You really have to sit back and ask yourself this question, how can anyone vote for Hillary, she lies to you, she lies about"
_blaairee|WeekendSchemers|-0.3818|0.245|0.755|0.0|RT @WeekendSchemers: This is embarrassing. Hillary vs Hillary https://t.co/59K9hRKTe7
_blaairee|twitter|-0.3818|0.245|0.755|0.0|RT @WeekendSchemers: This is embarrassing. Hillary vs Hillary https://t.co/59K9hRKTe7
DnbglrDian|KeithOlbermann|-0.6705|0.31|0.69|0.0|"RT @KeithOlbermann: Today's presidential ballot: Hillary Clinton, or national suicide: https://t.co/uBPp5vragL"
DnbglrDian|twitter|-0.6705|0.31|0.69|0.0|"RT @KeithOlbermann: Today's presidential ballot: Hillary Clinton, or national suicide: https://t.co/uBPp5vragL"
KarmaDrakpa|twitter|0.0|0.0|1.0|0.0|Translation:Question: Does Hillary wear red because shes a communist? #ElectionNight https://t.co/eFs3QJX41L
JaakeSweeney|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
JaakeSweeney|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
CarimarcelxA|vickto_willy|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
CarimarcelxA|t|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
Rachel_axl|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Rachel_axl|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
bonniebethdail3|DonaldTrumpNewz|-0.3182|0.228|0.642|0.13|"RT @DonaldTrumpNewz: Colin Powell TRUTH Revealed In Last Moments, Hillary Used Obama To HIDE Her Treason https://t.co/ZDWDfSazUK https://t."
bonniebethdail3|endingthefed|-0.3182|0.228|0.642|0.13|"RT @DonaldTrumpNewz: Colin Powell TRUTH Revealed In Last Moments, Hillary Used Obama To HIDE Her Treason https://t.co/ZDWDfSazUK https://t."
ALANLITTLE9|chadsdaddy|0.0|0.0|1.0|0.0|"RT @chadsdaddy: Savannah, Ga._Son just called VOTED TRUMP @noon today_checked ballot_switched to CROOKED HILLARY again on 2nd. attempt_ htt"
Tommy_Tsunami13|KayzoMusic|0.765|0.0|0.68|0.32|RT @KayzoMusic: If Hillary Clinton wins I hope she comes out for her victory speech to jotaro.
CarinaNicole16|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
CarinaNicole16|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
dracha|FrankLuntz|0.6369|0.0|0.733|0.267|"RT @FrankLuntz: The numbers I'm getting now suggest a nationwide turnout that strongly favors Hillary.And if Hillary does well, so will d"
Toddwagner14|Sam_Fridley14|-0.1695|0.074|0.926|0.0|"RT @Sam_Fridley14: ""The reason I voted for Hillary Clinton is because she is a woman."" This is not okay. This is not a legitimate reason."
inhalekidrauhl_|TheOneandOnIyUS|0.7096|0.0|0.753|0.247|RT @TheOneandOnIyUS: The joke is on Hillary if she wins. She'll have to sit at the desk Monica sat under.
Carrieecheungg|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
zzoerrose|AlexPisanti|-0.4404|0.153|0.847|0.0|RT @AlexPisanti: I'm scared I'm going to wake up and Hillary is going to be president #TrumpPence16
saucy_chica|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
_longdarrell|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
MichaelMcGan|DrMartyFox|-0.296|0.121|0.879|0.0|RT @DrMartyFox: #ImVotingBecause We Must Stop DUAL #JUSTICEWhere #Deplorables Must Follow The #RuleOfLawWhile #Hillary &amp; Her Cronies
Where_To_Now_|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Where_To_Now_|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
paully62|ananavarro|0.9351|0.0|0.496|0.504|@ananavarro Sweet Justice? And Hillary is such a good example and so inspiring and inclusive we should vote for her. Please.
Partywhatparty|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
UndyingCunt|BroHumors|0.0|0.0|1.0|0.0|ScreamingRT @BroHumors: Trump vs. Hillary  https://t.co/oVeD6xWBxL
UndyingCunt|vine|0.0|0.0|1.0|0.0|ScreamingRT @BroHumors: Trump vs. Hillary  https://t.co/oVeD6xWBxL
WareButch|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
arodgersw|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
arodgersw|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
vulnicore|OhNoSheTwitnt|0.4168|0.0|0.883|0.117|RT @OhNoSheTwitnt: Out to dinner in North Carolina wearing my Hillary shirt. It's under a sweater though I'm not stupid these people have g
AnnPettifor|Fullcarry|0.0772|0.0|0.874|0.126|RT @Fullcarry: Merkel May Yellen Hillary.... is that a proper sentence?
emilyb77|Hardline_Stance|0.6486|0.0|0.806|0.194|RT @Hardline_Stance: if Hillary wins not only will the BORDERS will be WIDE OPEN but she'll send letters all over the world inviting them o
bxnitvvpplebum_|RH1_ERA|0.5994|0.0|0.755|0.245|RT @RH1_ERA: How y'all voting for Bernie and Bernie voting for Hillary.. Lmao
vachilly64|dbk515|0.3818|0.0|0.847|0.153|RT @dbk515: Go Vote TodayLike for Hillary RT for Trump Please vote so we can get a big poll number #ElectionDay #Election2016 #Vote20
jpognon12|JerryGomezLope1|0.0|0.0|1.0|0.0|@JerryGomezLope1 Hillary Clinton
ludylugo|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
AndrewRR92|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
HarrisonCbryan|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
HarrisonCbryan|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Islandmike13|pablorodas|0.8436|0.0|0.702|0.298|RT @pablorodas: Hillary winning in 7 key states followed by Slate tracker! Great! #tcot #PJNET #GOP #2A #ccot #teaparty #tlot #MAGA #Trump2
majiktinkerbell|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @MaddieAndMichi @enjoynChi @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE
drgreenface|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
wolfiemouse|DeeStonewall|0.0|0.0|1.0|0.0|RT @DeeStonewall: #Bernie says #StrongerTogether#WeAreWithHer #Election2016 #Hillary#ClintonKaine2016 https://t.co/UoIMVkAgUR
wolfiemouse|twitter|0.0|0.0|1.0|0.0|RT @DeeStonewall: #Bernie says #StrongerTogether#WeAreWithHer #Election2016 #Hillary#ClintonKaine2016 https://t.co/UoIMVkAgUR
rihfashion|PopCrave|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
rihfashion|twitter|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
BradleyWasson|DrMartyFox|-0.3612|0.189|0.683|0.129|RT @DrMartyFox: #ImVotingBecause We Must Save Babies From #Hillary &amp; #PlannedParenthood Who Will Kill A Baby Minutes Before Birth &amp; S
MatiasAlegria3|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
MatiasAlegria3|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Spicoli83|megynkelly|0.0|0.0|1.0|0.0|@megynkelly rooting for Hillary @FoxNews She's past her prime #FireMegynKelly
FreedomTribe15|FredZeppelin12|0.4404|0.0|0.884|0.116|"RT @FredZeppelin12: This needs to be RT'dHillary Clinton: ""We're Going to Take Things Away From You on Behalf of the Common Good"" http:"
Johanna_Bowman|BernersUnited|0.5499|0.0|0.876|0.124|RT @BernersUnited: In my family 3 of us voted Stein and 1 voted for Hillary. We live in NY. NY always goes blue but hopefully stein will ge
kyle_blackman|YoungDems4Trump|0.0|0.0|1.0|0.0|RT @YoungDems4Trump: A message to both Democrats and Republicans:Voting against Hillary will be the most patriotic thing you'll ever do i
JoshNoneYaBiz|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
JoshNoneYaBiz|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
alohasusvn|jiujiuyulin|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
alohasusvn|twitter|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
Raheemc_|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Raheemc_|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
lufansloveluhan|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
crowjane29|pastemagazine|0.34|0.0|0.862|0.138|"Samantha Bee Endorses Hillary, Reads Emails and Goes to Russia In Last Pre-Election Full Frontal https://t.co/NXaTAibi8G"
americanyogini|isaacmojo|0.5984|0.0|0.72|0.28|@isaacmojo @Republiicunts @CorrectRecord I'm working with Hillary because she's a fucking hero.
amazinmind|amazinmind|0.4574|0.0|0.8|0.2|RT @amazinmind: Let's Go Nevada! Help Catherine give Hillary a Blue Senate majority. https://t.co/ALNbHNV5tu
amazinmind|twitter|0.4574|0.0|0.8|0.2|RT @amazinmind: Let's Go Nevada! Help Catherine give Hillary a Blue Senate majority. https://t.co/ALNbHNV5tu
TabacosCA|TabacosCA|-0.9317|0.517|0.483|0.0|RT @TabacosCA: HUMILIATION: HILLARY CAMP FREAKS OVER SHOCK PHOTO FROM CAMPAIGN RALLY SHOWING TOTAL FAILURE   https://t.co/9DwJm5NuEy https:
TabacosCA|youtube|-0.9317|0.517|0.483|0.0|RT @TabacosCA: HUMILIATION: HILLARY CAMP FREAKS OVER SHOCK PHOTO FROM CAMPAIGN RALLY SHOWING TOTAL FAILURE   https://t.co/9DwJm5NuEy https:
1johnfive|larryelder|0.6597|0.0|0.707|0.293|"RT @larryelder: In Other News: ""Grand Dragon Of California Of The KKK Endorses Hillary Clinton""https://t.co/NOzIMj6oMD#AnybodyButClinton"
1johnfive|usnews|0.6597|0.0|0.707|0.293|"RT @larryelder: In Other News: ""Grand Dragon Of California Of The KKK Endorses Hillary Clinton""https://t.co/NOzIMj6oMD#AnybodyButClinton"
amishabarnes2|chungaah|0.3818|0.122|0.667|0.211|RT @chungaah: Not even worried about the election Ik who gonna win Hillary obviously 
ArchangelMagicx|ObviousTwoll|-0.4019|0.137|0.863|0.0|"RT @ObviousTwoll: @RealJamesWoods not once has a ""calibration error"" turned a Hillary vote into a Trump vote. Soros resorting to desperatel"
ohmyzan|hyunascult|-0.5214|0.2|0.698|0.103|"@hyunascult like this entire election, even when BERNIE was running, she was all for Hillary so wtf is this"
bettyssd|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Obama continues Election Day ritual for Hillary Clinton https://t.co/uxU8EZ7jC3
bettyssd|washingtonpost|0.0|0.0|1.0|0.0|RT @washingtonpost: Obama continues Election Day ritual for Hillary Clinton https://t.co/uxU8EZ7jC3
kuhar_l|bfraser747|-0.7351|0.279|0.721|0.0|RT @bfraser747:  #NotAboveTheLaw #FBI agents are furious #Hillary wasn't indictment Director Comey has made #FBI look ridiculous #V
dabbinkook|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
cybranded|Bangelnuts|0.0|0.0|1.0|0.0|RT @Bangelnuts: #StayInLine Rock the vote for Hillary by staying in line.
spalienaceship|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
spalienaceship|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
Danielpm74|theScore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
Danielpm74|thescore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
xlarrykissx|csydelko|0.7506|0.0|0.758|0.242|RT @csydelko: 4 years ago I was on CNN for Obama's reelection. Hopefully I'll be making the same face when Hillary wins tonight. https://t.
xlarrykissx||0.7506|0.0|0.758|0.242|RT @csydelko: 4 years ago I was on CNN for Obama's reelection. Hopefully I'll be making the same face when Hillary wins tonight. https://t.
Cilveeuh_|twitter|0.0|0.0|1.0|0.0|I'm voting for Hillary because she pushed her  https://t.co/mFDa1SilM3
MeganOfTheOpera|FIirtationship|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
MeganOfTheOpera|twitter|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
DuesEmily|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
DuesEmily|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
jocemtzz|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
sirdrano|HaskelBiz|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
sirdrano|twitter|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
Gycez|YbsLucky|-0.8441|0.269|0.731|0.0|RT @YbsLucky: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
andrea_blake19|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
AnalissaVela|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
cats_executive|yankeebrit77|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
cats_executive|twitter|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
starwalker2012|thetruthdivision|-0.6523|0.348|0.652|0.0|EXIT POLL SHOCKER: Trump Beating Hillary By Incredible Margins In Florida https://t.co/R3ipxzGkm2
maaamoo_|TheAfghanDrake|-0.7121|0.229|0.771|0.0|RT @TheAfghanDrake: Vote for Hillary Clinton. I don't care if she's a liar or sketchy. Y'all boyfriends lie to y'all everyday and y'all sti
camhoops1|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
amigoalfil|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: ""If you believe we should never write discrimination into our laws...youve got to vote! Hillary https://t.co/jfd3CXL"
amigoalfil|t|0.0|0.0|1.0|0.0|"RT @HillaryClinton: ""If you believe we should never write discrimination into our laws...youve got to vote! Hillary https://t.co/jfd3CXL"
karindarby|DineshDSouza|0.0|0.0|1.0|0.0|"RT @DineshDSouza: IT'S UP TO US: We can't rely on others to do our work; we have to do our work--on Tuesday, the American people are Hillar"
kelsey_ryan20|SirGabrielofLO|0.857|0.0|0.692|0.308|RT @SirGabrielofLO: Will Hillary win by a landslide? Can Trump make American great again? Netflix ever have updated movies? Find out next t
miflorhermosa|SInow|0.0|0.0|1.0|0.0|RT @SInow: Colin Kaepernick said he isnt voting in the election https://t.co/9IfZWrKNCc https://t.co/l3kO9BORir
miflorhermosa|si|0.0|0.0|1.0|0.0|RT @SInow: Colin Kaepernick said he isnt voting in the election https://t.co/9IfZWrKNCc https://t.co/l3kO9BORir
AMWG9|laurenasarson|-0.6022|0.275|0.595|0.129|"@laurenasarson Most people care more about actions instead of words. Trumps words were bad, Hillary left 4 people to die."
BellaLucky4|Pamela_Moore13|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
BellaLucky4|twitter|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
televisedprogrm|triciavicious|0.5719|0.0|0.709|0.291|RT @triciavicious: if Hillary wins I'm leaking my own nudes
oriori1697|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
oriori1697|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
RiverRatWA57|twitter|0.0|0.0|1.0|0.0|VOTE TRUMP VOTE TRUMP VOTE TRUMP VOTE TRUMP NOW!!!!!!!!!!!!Hillary for Prison!!!!! https://t.co/lQAY7ZIlZs
ansguevarra1|CoreyGrossJr|0.7955|0.0|0.56|0.44|@CoreyGrossJr Whoever who wins it's under God's hands.. Hoping Hillary !!
MoneyMills_72|ashleysharpen|0.0772|0.0|0.902|0.098|RT @ashleysharpen: It blows my mind that people actually want Hillary in office
carolinekjones|TheDonaldNews|0.0|0.0|1.0|0.0|RT @TheDonaldNews: KENTUCKY : 68% TRUMP ------ 28% HILLARY https://t.co/ERKVVnh1PL
carolinekjones|twitter|0.0|0.0|1.0|0.0|RT @TheDonaldNews: KENTUCKY : 68% TRUMP ------ 28% HILLARY https://t.co/ERKVVnh1PL
PantsuitEnFuego|theothermurph51|-0.8156|0.364|0.582|0.054|"RT @theothermurph51: @RawStory Hey @MichelleObama , that's the point!We arent playing round! We want #Hillary 2 lose &amp; go 2 prison!!"
jetblacklovato|vibeeeez|-0.5574|0.261|0.739|0.0|RT @vibeeeez: prediction: Hillary Clinton is our next present &amp; everyone is shocked Trump lost
DrThomasPaul|DrThomasPaul|0.0|0.0|1.0|0.0|RT @DrThomasPaul: All that the uniformed have are projections of unresolved issues which belong in #THERAPY sessions. #Hillary #Trump https
Mrgee_bande|JOHNSONSFOOL|0.7579|0.0|0.727|0.273|"RT @JOHNSONSFOOL: you still have time, please please go vote for hillary, she's the better option for you &amp; the youths future #ElectionNigh"
r1965rainey|gdweo|0.0|0.0|1.0|0.0|RT @gdweo: Drove 700 miles to get your vote in-Lots of ppl won't even walk to the end of the driveway-Those deserve a Hillary America https
nochillvalerie|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
nochillvalerie|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
RobertMabr|JustMe3316|0.0|0.0|1.0|0.0|@JustMe3316 @MiceeMouse @JimPowersjpp @thegreatfeather  @Promo_Bob_ the hillary wrap has been known to burst into flames even in a rainstorm
starknightz|foxnews|0.0|0.0|1.0|0.0|BREAKING! POLL LOCKDOWN IN S. California after shooting https://t.co/s8rv1bKuf4 #hillary #Trump #ElectionNight #TrumpTrain
Iocalwhiteboy|britishdcddy|0.0|0.0|1.0|0.0|@britishdcddy I rooting for Hillary in reality. But I did bet $5 on trump just because.
ashxbandz|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
ashxbandz|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
PeriodicaI|nytimes|0.0|0.0|1.0|0.0|How the FBI Reviewed Thousands of Emails in One Week - New York Times https://t.co/xmF5IkAP95
samavsfan|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
samavsfan|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
scifical|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
scifical|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
saragomezzzz|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
HmrncnrnHolli|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
happykt|FelicityHuffman|0.7371|0.0|0.633|0.367|RT @FelicityHuffman: Voter loveWE LOVE HILLARY! @HillaryClinton #electionday #ImWithHer https://t.co/0AaJTaubSe
happykt|twitter|0.7371|0.0|0.633|0.367|RT @FelicityHuffman: Voter loveWE LOVE HILLARY! @HillaryClinton #electionday #ImWithHer https://t.co/0AaJTaubSe
auztinphillips|TheWizKhalifa|-0.9022|0.41|0.59|0.0|RT @TheWizKhalifa: People hate Trump because the media made them hate Trump.People hate Hillary because they are paying attention.#Elec
garbagecuntt|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
DanielOzioma6|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
DanielOzioma6|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
GutsyJupiter49|AltStreamMedia|-0.2787|0.172|0.661|0.167|"RT @AltStreamMedia: #ImVotingBecause they can't. Stop Hillary, stop war. Rebuild our country at home. Let's do this. https://t.co/xDH4Nin1cu"
GutsyJupiter49|twitter|-0.2787|0.172|0.661|0.167|"RT @AltStreamMedia: #ImVotingBecause they can't. Stop Hillary, stop war. Rebuild our country at home. Let's do this. https://t.co/xDH4Nin1cu"
usvoteout|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana: 0.9% reporting TRUMP 70.5% | Hillary 25.8% massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Elect
PrynxRex|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
HRC1947|lizcgoodwin|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
HRC1947|twitter|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
DaphneBinulski|RepCoriFournier|0.0|0.0|1.0|0.0|RT @RepCoriFournier: This is what @CNN is counting on with the BIG push on their network that Republicans will be voting HILLARY n republic
xileenie|ppetrov5|0.0|0.0|1.0|0.0|"RT @ppetrov5: Hillary Clinton and her campaign met with prioritiesUSA, which is against the law. #PodestaEmails35 #wikileaks #fbi https://t"
xileenie||0.0|0.0|1.0|0.0|"RT @ppetrov5: Hillary Clinton and her campaign met with prioritiesUSA, which is against the law. #PodestaEmails35 #wikileaks #fbi https://t"
Mikmunt|Pudingtane|0.0|0.0|1.0|0.0|RT @Pudingtane: BREAKING-hillary-clintons-$20-million-0bama-bribe-to-become-us-secretary-of-state-leaked-by-fbi. https://t.co/7v7kiPCD7n
Mikmunt|endingthefed|0.0|0.0|1.0|0.0|RT @Pudingtane: BREAKING-hillary-clintons-$20-million-0bama-bribe-to-become-us-secretary-of-state-leaked-by-fbi. https://t.co/7v7kiPCD7n
QGS24|joe_fortkort5|0.1655|0.089|0.759|0.152|RT @joe_fortkort5: People love to talk about Hillary and Trump and how important this election is but forget the Warriors blew a 3-1 lead i
squidninja|healthandcents|0.3885|0.186|0.522|0.292|RT @healthandcents: #ElectionFinalThoughtsI #ImVotingBecause Hillary LET FOUR HEROES DIE #Benghazi POTUS #Trump SUPPORTS #Military &amp; #V
hillary_gibble|mdj17|0.0|0.0|1.0|0.0|"RT @mdj17: Government Workers Now Outnumber Manufacturing Workers by 9,977,000THE SIGN WE ARE APPROACHING SOCIALISM  https://t.co/2R3EA8O"
hillary_gibble|t|0.0|0.0|1.0|0.0|"RT @mdj17: Government Workers Now Outnumber Manufacturing Workers by 9,977,000THE SIGN WE ARE APPROACHING SOCIALISM  https://t.co/2R3EA8O"
phichitxt|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
NewSonOfLiberty|newsmax|0.0|0.0|1.0|0.0|"RT @newsmax: With 1% of the vote in for Kentucky, Trump is holding a steady lead over Hillary Clinton. #ElectionNight #myvote2016 https://t"
NewSonOfLiberty||0.0|0.0|1.0|0.0|"RT @newsmax: With 1% of the vote in for Kentucky, Trump is holding a steady lead over Hillary Clinton. #ElectionNight #myvote2016 https://t"
YoungMooo|_iAmRoyal|-0.8957|0.329|0.671|0.0|"RT @_iAmRoyal: Right now, Hillary is threatening to go to war with several countries. She's JUST as bad as Trump depending on who you ask."
ToplessGoddess|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
ToplessGoddess|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
donnalea1788|Lrihendry|0.7256|0.0|0.738|0.262|"RT @Lrihendry: Hillary supports this! If this is reason enough to support Trump, then you might want to sit this one out! #ElectionFina"
Maine4Trump|kincannon_show|-0.5849|0.296|0.704|0.0|RT @kincannon_show: This is very bad for Hillary --&gt; https://t.co/lv5ybXLiHZ
Maine4Trump|twitter|-0.5849|0.296|0.704|0.0|RT @kincannon_show: This is very bad for Hillary --&gt; https://t.co/lv5ybXLiHZ
jazlynrxzo|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
OCEANGRIMEZ|notmily|-0.1531|0.133|0.719|0.147|RT @notmily: i hate donald trump and hillary clinton we are better off all going back to england and apologising for what we've done
_marsh_y|drefamous|-0.1027|0.06|0.94|0.0|RT @drefamous: if Rihanna wearing a shirt with Rihanna wearing a shirt with Hillary Clinton on it doesnt make ur day then idk what will. h
_JasonAA|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
butleriano|jiujiuyulin|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
butleriano|twitter|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
froggyboyfriend|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
manicsocratic|theslot|-0.7269|0.357|0.643|0.0|"All the Sad, Woke Men Forced to Vote for Hillary Clinton https://t.co/fRP4VrrMgm https://t.co/yWjTFGeB85"
TheSolClarke|ameeritalsham|-0.4215|0.138|0.804|0.058|"RT @ameeritalsham: Hillary Clinton: ""I want the Iranians to know, that if I'm the president, we will attack Iran"" https://t.co/FMb2jIqIRF"
TheSolClarke|twitter|-0.4215|0.138|0.804|0.058|"RT @ameeritalsham: Hillary Clinton: ""I want the Iranians to know, that if I'm the president, we will attack Iran"" https://t.co/FMb2jIqIRF"
Benhur_Gill|realDonaldTrump|0.0|0.0|1.0|0.0|Come on #Utah@realDonaldTrump needs every single last vote!We cannot let Hillary have UtahIt may begin &amp; end wit https://t.co/hpU11pqnzE
Benhur_Gill|twitter|0.0|0.0|1.0|0.0|Come on #Utah@realDonaldTrump needs every single last vote!We cannot let Hillary have UtahIt may begin &amp; end wit https://t.co/hpU11pqnzE
jamieraegomes|dezlsmith|0.7184|0.0|0.684|0.316|RT @dezlsmith: Voted and pray Hillary wins. Trump Presidency is a nightmare we won't survive  #ElectionNight
Hals115|hyatt_jonathan|-0.4449|0.197|0.803|0.0|RT @hyatt_jonathan: If Hillary couldn't even please Bill what makes anybody believe she could please our county? #Hillary4Prison
jadawarren13|StevannaA|0.3832|0.101|0.71|0.189|RT @StevannaA: It blows my mind that so many Americans who were raised to value honesty are completely ignoring the fact that Hillary CANNO
PeriodicaI|usatoday|0.197|0.0|0.861|0.139|Hillary Clinton calls voting for herself a 'most humbling feeling' - USA TODAY https://t.co/H70Ojke1Ob
JMonet__|MannequinVid|0.0|0.0|1.0|0.0|RT @MannequinVid: Hillary Clinton #MannequinChallenge  https://t.co/9ipPwXdqEi
JMonet__|twitter|0.0|0.0|1.0|0.0|RT @MannequinVid: Hillary Clinton #MannequinChallenge  https://t.co/9ipPwXdqEi
kori_martez|___DestinyJadai|-0.6739|0.476|0.524|0.0|"RT @___DestinyJadai: ""VOTE HILLARY BITCH""  https://t.co/xVltWc6dU7"
kori_martez|twitter|-0.6739|0.476|0.524|0.0|"RT @___DestinyJadai: ""VOTE HILLARY BITCH""  https://t.co/xVltWc6dU7"
SeanFleming1916|ltsDonaIdTrump_|0.0|0.0|1.0|0.0|RT @ltsDonaIdTrump_: Hillary Clinton's da sells avon
antionettemat10|twitter|0.0|0.0|1.0|0.0|Me too..gooooooooooo Hillary https://t.co/uVGwZKf07a
mamasaurusof2|MMFlint|-0.4019|0.119|0.881|0.0|RT @MMFlint: The word throughout Michigan has been long lines in Hillary neighborhoods and long lines in the deer blind hoods.
DanielChappers|SoVeryFinnish|0.4019|0.0|0.787|0.213|RT @SoVeryFinnish: When you live in Nurmijrvi and support Hillary. https://t.co/878erqvj8M
DanielChappers|twitter|0.4019|0.0|0.787|0.213|RT @SoVeryFinnish: When you live in Nurmijrvi and support Hillary. https://t.co/878erqvj8M
iStayClassyOH|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
iStayClassyOH|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Mr3lsewhere|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Mr3lsewhere|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
AndrewsCosta4|TheSun|0.6204|0.0|0.807|0.193|RT @TheSun: A final poll for the #USElection shows who is most likely to win tonight #USElection https://t.co/6cWAQBvrhi https://t.co/AchWa
AndrewsCosta4|thesun|0.6204|0.0|0.807|0.193|RT @TheSun: A final poll for the #USElection shows who is most likely to win tonight #USElection https://t.co/6cWAQBvrhi https://t.co/AchWa
da11asc|twitter|0.0|0.0|1.0|0.0|you already chose hillary  https://t.co/MZ583CWSzO
__lizbethxo|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
__lizbethxo|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
HarmoHeather|LindforLind|-0.4767|0.119|0.881|0.0|RT @LindforLind: To me it's not a big deal that Hillary is a woman. The big deal is that Donald Trump is toxic and dangerous. #ElectionNight
savannahsand3rs|twitter|-0.5859|0.655|0.345|0.0|wtf Hillary https://t.co/s5AiQRbDQ3
magssnider|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
NotoriousMNR|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
NotoriousMNR|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
BeySickening|beyupdates_|0.3612|0.0|0.815|0.185|RT @beyupdates_: Me: *votes for Hillary* Hillary: Thank you for vot-Me: https://t.co/nx99GlD5gc
BeySickening|twitter|0.3612|0.0|0.815|0.185|RT @beyupdates_: Me: *votes for Hillary* Hillary: Thank you for vot-Me: https://t.co/nx99GlD5gc
Y0SHIHARA|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Y0SHIHARA|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ouhshejocelyn|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
MamiPerkins|vickto_willy|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
MamiPerkins|t|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
SHaMRecKs|FFrantec|0.4404|0.221|0.41|0.369|@FFrantec @zThumperr hillary is a whore she guzzles cum for fun lmao
wendtoverthere|twitter|0.0|0.0|1.0|0.0|"""I'm voting for Trump because he's not Hillary""""I'm voting for Hillary because she's not Trump"" https://t.co/M0YPfjzzrT"
kylieslipkit|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
kylieslipkit|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Austin_Gilstrap|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Austin_Gilstrap|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
BillKS1|umpire43|0.0|0.0|1.0|0.0|RT @umpire43: A woman in Fla reported she voted Trump on Smartmatic https://t.co/Sm6mmsb0AH was flipped to Hillary and multiplied to 200 in
BillKS1||0.0|0.0|1.0|0.0|RT @umpire43: A woman in Fla reported she voted Trump on Smartmatic https://t.co/Sm6mmsb0AH was flipped to Hillary and multiplied to 200 in
elaine_wildes|asdomke|-0.6249|0.282|0.718|0.0|RT @asdomke: Polls disappear showing major Hillary collapse among likely voters on election day... https://t.co/zI3JeNYMCO
elaine_wildes|linkis|-0.6249|0.282|0.718|0.0|RT @asdomke: Polls disappear showing major Hillary collapse among likely voters on election day... https://t.co/zI3JeNYMCO
le_american|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
le_american|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
Baxenwald|ppyajunebug|-0.2244|0.136|0.864|0.0|RT @ppyajunebug: 2016Trump: No man but I can lead this country to greatness!Hillary: https://t.co/EINQIRMg8o
Baxenwald|twitter|-0.2244|0.136|0.864|0.0|RT @ppyajunebug: 2016Trump: No man but I can lead this country to greatness!Hillary: https://t.co/EINQIRMg8o
byrnesmaeve06|sassytbh|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
byrnesmaeve06|twitter|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
dmshea|THR|0.7003|0.0|0.674|0.326|RT @THR: #ElectionDay: Hillary Clinton thanks Facebook supporters known as the #PantsuitNation https://t.co/imJyIz3QPM https://t.co/xMnObze
dmshea|hollywoodreporter|0.7003|0.0|0.674|0.326|RT @THR: #ElectionDay: Hillary Clinton thanks Facebook supporters known as the #PantsuitNation https://t.co/imJyIz3QPM https://t.co/xMnObze
laurendorwart|CloydRivers|0.0|0.0|1.0|0.0|RT @CloydRivers: Im not against a woman bein President. Im just against that woman bein Hillary Clinton. Merica.
lezmone|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
CubsFanJohn|CNNPolitics|0.0|0.0|1.0|0.0|"RT @CNNPolitics: George W. Bush did not vote for Clinton, despite what Rush Limbuagh claims https://t.co/5FhnosgEh4 https://t.co/vOvJQZEUxA"
CubsFanJohn|money|0.0|0.0|1.0|0.0|"RT @CNNPolitics: George W. Bush did not vote for Clinton, despite what Rush Limbuagh claims https://t.co/5FhnosgEh4 https://t.co/vOvJQZEUxA"
MackCollier|CNN|0.0|0.0|1.0|0.0|".@CNN will start calling states immediately for Hillary in a few mins.  Bogus, your vote counts esp in Mountain &amp; West Coast #electionnight"
1975jetsfan4|twitter|0.8294|0.0|0.571|0.429|"Okay for LeBron &amp; Hollywood supporting Hillary but not for Belichick to support Trump?  Ok, hypocrite. https://t.co/6yYBsgeFy9"
hopelmez16|dougsmith1946|0.0|0.0|1.0|0.0|RT @dougsmith1946: @nationdivided @janiehburton  @FBI @FBIWFO  @NewYorkFBI  That's why officials stuffed ballot boxes for Hillary https://t
hopelmez16||0.0|0.0|1.0|0.0|RT @dougsmith1946: @nationdivided @janiehburton  @FBI @FBIWFO  @NewYorkFBI  That's why officials stuffed ballot boxes for Hillary https://t
jetblacklovato|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
jetblacklovato|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
ally_gardener|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
JohnTrumpFanKJV|mitchellvii|-0.3182|0.206|0.653|0.141|"RT @mitchellvii: If true, this is brutal for Hillary.  She won't match Obama's numbers. https://t.co/z0o069Bv1p"
JohnTrumpFanKJV|twitter|-0.3182|0.206|0.653|0.141|"RT @mitchellvii: If true, this is brutal for Hillary.  She won't match Obama's numbers. https://t.co/z0o069Bv1p"
notbuyingthat54|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
rachelevans_28|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
AndresUseche|Digg|-0.1531|0.082|0.918|0.0|Pregnant woman votes 4 #Hillary while in labour after stopping at polls en route to hospital #electionday https://t.co/7ZBqblt2bx via @Digg
AndresUseche|telegraph|-0.1531|0.082|0.918|0.0|Pregnant woman votes 4 #Hillary while in labour after stopping at polls en route to hospital #electionday https://t.co/7ZBqblt2bx via @Digg
__FinesseKvng|GIRLHEFUNNY|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
__FinesseKvng|twitter|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
rosegoggles|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
rosegoggles|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
anndddreaaa|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
CrossFit4PRO|Inc|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
CrossFit4PRO|t|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
leighsm84975411|NickOchsnerWBTV|0.5859|0.0|0.798|0.202|@NickOchsnerWBTV @WBTV_News yea just keep it open until you get enough votes for Hillary to win.
CrookedOrange|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
CrookedOrange|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
WamplerJim|BobMacAZ|-0.6908|0.239|0.761|0.0|"RT @BobMacAZ: BREAKING: Hours Before Polls Close, Rape Allegation Sends Hillary Into Tailspin https://t.co/sU3y6q2Bu7 via @USADailyInfo"
WamplerJim|dailyinfo|-0.6908|0.239|0.761|0.0|"RT @BobMacAZ: BREAKING: Hours Before Polls Close, Rape Allegation Sends Hillary Into Tailspin https://t.co/sU3y6q2Bu7 via @USADailyInfo"
yourBAD_habbit|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
tweetwithtee|WayneL_Jr|0.0|0.0|1.0|0.0|RT @WayneL_Jr: I think it's time to put her down RT @luke_santa: My grandma after someone vandalized her house w/ a Hillary sign https://t.
tweetwithtee||0.0|0.0|1.0|0.0|RT @WayneL_Jr: I think it's time to put her down RT @luke_santa: My grandma after someone vandalized her house w/ a Hillary sign https://t.
vylancex|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
vylancex|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
CrownMeTaylor|GIRLHEFUNNY|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
CrownMeTaylor|twitter|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
USAHipster|PrisonPlanet|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
USAHipster|pittsburgh|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
danihertz88|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
Diane401k|courierjournal|-0.6908|0.289|0.711|0.0|"RT @courierjournal: Joshua Roy, 18, said he's tired of all of Hillary's lies https://t.co/Ger1DjwX9n #KyElect #InElect"
Diane401k|courier-journal|-0.6908|0.289|0.711|0.0|"RT @courierjournal: Joshua Roy, 18, said he's tired of all of Hillary's lies https://t.co/Ger1DjwX9n #KyElect #InElect"
HadleyKiefer|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
HadleyKiefer|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
NECN|necn|0.0|0.0|1.0|0.0|WATCH LIVE: necn's election night coverage. https://t.co/TjMPutYNa0
OKC_luver_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
OKC_luver_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
caseyyy_h|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
caseyyy_h|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
BlackbirdHarm|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
efairhurst|money|0.0|0.0|1.0|0.0|"Hillary Clinton's mostly female press corps on covering 'big moment in history' - Nov. 8, 2016 https://t.co/5zobdU2kmJ"
SophieSwancott9|freckledbutt|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
SophieSwancott9|twitter|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
APettyQueen|facebook|-0.5023|0.244|0.641|0.114|"Hillary is not ""better"" than Trump. Trump is not some horrible guy because he's racist, sexist, ignorant and... https://t.co/EiE766BvpS"
707spookyboo22|verizon|0.3129|0.164|0.602|0.234|@verizon oh look! it's the map that is going to defeat hillary! yay!
casey2513|ReturnofRV|0.1779|0.109|0.746|0.144|"RT @ReturnofRV: Why are all the Hillary supporters, Hillary trolls, and Hillary mainstream media pundits strangely quiet?"
corruptvoltaire|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
Keithmadigan|billmaher|-0.8753|0.382|0.574|0.044|"RT @billmaher: Pls vote for Hillary today. Even if you don't like her, its necessary to block a dangerous lunatic ultimate power. #ThisTime"
TrlnWatermelon|pops_clark|0.765|0.0|0.664|0.336|RT @pops_clark: @darkagesreturn Thanks. Wifey fine. Right now exit polls show slaughter. 83%Trump. 13% Hillary. Looks real good.
john_bugaj|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
biebstorture|jaureologist|-0.0516|0.207|0.591|0.202|RT @jaureologist: I DON'T CARE HOW MUCH Y'ALL HATE BOTH CANDIDATES YOU WILL VOTE FOR HILLARY WHETHER YOU LIKE IT OR NOT I REFUSE TO LET TRU
frespirit01|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @YoungDems4Trump @enjoynChi @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE
TheWeek|theweek|0.6808|0.0|0.616|0.384|Hillary Clinton has a special message for her Pantsuit Nation supporters: https://t.co/UQb5tOq5zx
Yajasaher|mitchellvii|0.6597|0.0|0.735|0.265|"RT @mitchellvii: How can anyone think of trainwreck Hillary as a ""strong Commander in Chief""?  I mean, my God."
JoshNoneYaBiz|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
JoshNoneYaBiz|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
cloudydino|KayzoMusic|0.765|0.0|0.68|0.32|RT @KayzoMusic: If Hillary Clinton wins I hope she comes out for her victory speech to jotaro.
ButteryyToast|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
keith_camic|TeamTrump|0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
keith_camic||0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
ButerasThief|_actually_ash|-0.8402|0.267|0.733|0.0|@_actually_ash I'm for trump but this is a bad argument because at the time Hillary was a lawyer it was her job to cover it up
douglasnotdoug|bruner_sara4|0.9246|0.0|0.573|0.427|"RT @bruner_sara4: definitely rooting for hillary, but i think it's pretty important if she wins to not overlook her flaws/why people are so"
LindsayrenzLr|lizcgoodwin|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
LindsayrenzLr|twitter|0.0|0.0|1.0|0.0|"RT @lizcgoodwin: Hillary Clinton left a message to the women of the ""pantsuit nation"" Facebook group https://t.co/1CGPiX6BO3"
MimiieLafayette|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
MimiieLafayette|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
sag2horses|US_Army_Vet|0.0|0.0|1.0|0.0|RT @US_Army_Vet: Hillary had her maid print classified mat'l: NYPhttps://t.co/lEur7MncMo Breitbarthttps://t.co/q2nerd6kVU @American1765 @
marisawhittt|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
differentalexis|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
JohnCzer1|ldbrillante|0.5837|0.0|0.859|0.141|RT @ldbrillante: Hillary &amp; Trump are friend &amp; connected. You can't get rid of one by voting for the other!Reject the SCAM!Vote Dr. Jill S
_laurennewsome|ltsDonaIdTrump_|0.0|0.0|1.0|0.0|RT @ltsDonaIdTrump_: Hillary Clinton's da sells avon
MesutOzilexis|EmanDaGoon|-0.6597|0.386|0.614|0.0|RT @EmanDaGoon: Trump or Hillary. You're fucked America 
RubenHolguin29|instagram|0.5719|0.0|0.764|0.236|History will be made once again today when Hillary Clinton Wins as https://t.co/tXqsFPaBRk
ResetPolitics|BDUTT|0.4019|0.0|0.886|0.114|RT @BDUTT: Live from the Glass Ceiling I bet Hillary Clinton Will Smash tonight. The venue of her Victory Party. Facebook Live https://t.co
ResetPolitics|t|0.4019|0.0|0.886|0.114|RT @BDUTT: Live from the Glass Ceiling I bet Hillary Clinton Will Smash tonight. The venue of her Victory Party. Facebook Live https://t.co
MiikeTasticle|Soulovillain|-0.5994|0.163|0.837|0.0|RT @Soulovillain: She need to die already. RT @luke_santa My grandma's reaction after someone vandalized her house with a Hillary sign http
chill_kbye|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
blondediamond99|HillaryforMO|0.7783|0.0|0.726|0.274|RT @HillaryforMO: A vote for Hillary and Democrats down the ballot is a vote for the values that make America great: https://t.co/mVMj1fCCf
blondediamond99|t|0.7783|0.0|0.726|0.274|RT @HillaryforMO: A vote for Hillary and Democrats down the ballot is a vote for the values that make America great: https://t.co/mVMj1fCCf
Future_Boone|byalexus_|0.0|0.0|1.0|0.0|RT @byalexus_: Hillary is the next president.
liyuanwei|qz|0.0|0.0|1.0|0.0|RT @qz: From Nina Simone to Beyonce: The Quartz playlist of songs by women who rule https://t.co/34y9D4BdxT
liyuanwei|qz|0.0|0.0|1.0|0.0|RT @qz: From Nina Simone to Beyonce: The Quartz playlist of songs by women who rule https://t.co/34y9D4BdxT
DrThomasPaul|DrThomasPaul|0.0|0.0|1.0|0.0|RT @DrThomasPaul: .@realDonaldTrump #Trump's the kind of guy who will take you to #battle if necessary and then make you his #ally. He's a
kf4bef|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
ilbznu3|twitter|0.0|0.0|1.0|0.0|we getit wegetit wegotit...neither hillary nor theTrumper https://t.co/BaVKqMbg4U
soteruh|twitter|0.0|0.0|1.0|0.0|#MyVote2016 Not Hillary  #MAGA https://t.co/gDNZDYYHYt
mikemavroulis|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
okayskip|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
okayskip|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
nwts1224|KyraLawrence2|0.6124|0.0|0.762|0.238|RT @KyraLawrence2: Well since Hillary ran for president this time i better be seeing Michelle Obama in four years .
TonyBeavers1|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
guuurrrrrddds|kimayad_|0.3612|0.0|0.872|0.128|"RT @kimayad_: Before Hillary Clinton, there was Shirley Chisholm. Thank you for paving the way. #UnboughtAndUnbossed72 #Election2016 http"
BillJohnson42|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
BillJohnson42|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
BlueSeaSailing|ObviousTwoll|-0.4019|0.137|0.863|0.0|"RT @ObviousTwoll: @RealJamesWoods not once has a ""calibration error"" turned a Hillary vote into a Trump vote. Soros resorting to desperatel"
arusso1984|LisaEdelstein|0.8541|0.0|0.645|0.355|@LisaEdelstein can I ask you a question? Who do you think will win between Hillary and Trump? Thanks for the answer :-)
Armandoayala13|Truthbytony|-0.5859|0.297|0.703|0.0|RT @Truthbytony: Today's the day bitch. VOTE FA HILLARY. https://t.co/JSlc6ZCFrU
Armandoayala13|twitter|-0.5859|0.297|0.703|0.0|RT @Truthbytony: Today's the day bitch. VOTE FA HILLARY. https://t.co/JSlc6ZCFrU
badIandwentz|csydelko|0.7506|0.0|0.758|0.242|RT @csydelko: 4 years ago I was on CNN for Obama's reelection. Hopefully I'll be making the same face when Hillary wins tonight. https://t.
badIandwentz||0.7506|0.0|0.758|0.242|RT @csydelko: 4 years ago I was on CNN for Obama's reelection. Hopefully I'll be making the same face when Hillary wins tonight. https://t.
PilotJonesss_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
PilotJonesss_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ExtremeFit4life|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
ExtremeFit4life|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
_kassidywright_|jessicas1540|0.3612|0.0|0.872|0.128|RT @jessicas1540: could never vote for hillary clinton just for the fact of how much she supports abortions
superbrian75|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
superbrian75|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
raphaellaN|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
raphaellaN|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
Enger1776|SophiaHelwani|0.6696|0.0|0.781|0.219|RT @SophiaHelwani: Hillary's greatest hits #7. Obama does the okie doke songl!  @placeboing @joerogan @TimKennedyMMA @Cowboycerrone @mitche
RichardDBK|RichardDBK|-0.2732|0.091|0.864|0.045|"@RichardDBK No matter what you think of Hillary, that should at least give you pause to think about how historic this election is."
LepsJack|iduitmann|0.5719|0.0|0.821|0.179|RT @iduitmann: joke's on Hillary if she wins. she'll have to sit at the desk Monica sat under.
kiuwalsh|courierjournal|-0.6908|0.289|0.711|0.0|"RT @courierjournal: Joshua Roy, 18, said he's tired of all of Hillary's lies https://t.co/Ger1DjwX9n #KyElect #InElect"
kiuwalsh|courier-journal|-0.6908|0.289|0.711|0.0|"RT @courierjournal: Joshua Roy, 18, said he's tired of all of Hillary's lies https://t.co/Ger1DjwX9n #KyElect #InElect"
reneegoldsbery|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
JoeSaferly|realDonaldTrump|-0.2695|0.162|0.725|0.113|RT @realDonaldTrump: Hey Missouri let's defeat Crooked Hillary &amp; @koster4missouri! Koster supports Obamacare &amp; amnesty! Vote outsider Navy
TinaJ4Trump|TheDonaldNews|0.0|0.0|1.0|0.0|RT @TheDonaldNews: NEW HAMPSHIRE : 52% TRUMP   -----   41% HILLARY https://t.co/xNpCXbnHuR
TinaJ4Trump|twitter|0.0|0.0|1.0|0.0|RT @TheDonaldNews: NEW HAMPSHIRE : 52% TRUMP   -----   41% HILLARY https://t.co/xNpCXbnHuR
daiseyjane13|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
BobbyByThePound|Chubb_longway2|-0.5719|0.425|0.392|0.183|RT @Chubb_longway2: Trump is beating Hillary ass bro lol
Tweets_By_Zo|Jezebel|-0.7269|0.319|0.681|0.0|"RT @Jezebel: All the sad, woke men forced to vote for Hillary Clinton https://t.co/X22INC8Dqa https://t.co/LXAvCNzHX0"
Tweets_By_Zo|theslot|-0.7269|0.319|0.681|0.0|"RT @Jezebel: All the sad, woke men forced to vote for Hillary Clinton https://t.co/X22INC8Dqa https://t.co/LXAvCNzHX0"
Savageassnecy|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
Moviewatcher21|PrisonPlanet|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
Moviewatcher21|pittsburgh|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
weeeendyy_|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
weeeendyy_|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
RICindylou|stephenWalt|0.3612|0.0|0.8|0.2|@stephenWalt Probably be like his birther one. I concede to Hillary period.
ts65136|2ALAW|-0.5859|0.192|0.808|0.0|RT @2ALAW: Voter Fraud In PhiladelphiaPush Button One For HillaryPaid For By The Democratic County.#ElectionNight #DonaldTrump https:/
ts65136||-0.5859|0.192|0.808|0.0|RT @2ALAW: Voter Fraud In PhiladelphiaPush Button One For HillaryPaid For By The Democratic County.#ElectionNight #DonaldTrump https:/
mpanighetti|Spacekatgal|0.5106|0.0|0.875|0.125|"RT @Spacekatgal: CSPAN is passing out free copies of the constitution at Hillary HQ, which is the most C-SPAN thing to do ever. #ImWithHer"
lIbby_annn|MrDane1982|0.0|0.0|1.0|0.0|RT @MrDane1982: Niece: Uncle Dane I voted in pre school today for Hillary Clinton!! https://t.co/hGKpI0Fv8P
lIbby_annn|twitter|0.0|0.0|1.0|0.0|RT @MrDane1982: Niece: Uncle Dane I voted in pre school today for Hillary Clinton!! https://t.co/hGKpI0Fv8P
c38372346|MissLizzyNJ|0.0|0.0|1.0|0.0|RT @MissLizzyNJ: Oh so being married to a misogynistic serial adulterer makes Hillary a self-respecting woman? Give me a break. https:/
c38372346||0.0|0.0|1.0|0.0|RT @MissLizzyNJ: Oh so being married to a misogynistic serial adulterer makes Hillary a self-respecting woman? Give me a break. https:/
dejalenet|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
dejalenet|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
deessssst|pizzaparacenar|0.0|0.0|1.0|0.0|RT @pizzaparacenar: Ni Trump ni Hillary https://t.co/O4X2zybhAX
deessssst|twitter|0.0|0.0|1.0|0.0|RT @pizzaparacenar: Ni Trump ni Hillary https://t.co/O4X2zybhAX
dianuuhh|REALBrianStreng|0.7096|0.0|0.789|0.211|RT @REALBrianStreng: Joke is on Hillary if she wins the election because that means she has to sit at the desk Monica was under
styIesIuxe|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
RaylanWest|twitter|0.0|0.0|1.0|0.0|Hillary took money from Saudis. #WTFAmericaIn5Words https://t.co/0eNYVsHpkq
Laurie_LDL|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
Laurie_LDL|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
darthmiho|Spacekatgal|0.5106|0.0|0.875|0.125|"RT @Spacekatgal: CSPAN is passing out free copies of the constitution at Hillary HQ, which is the most C-SPAN thing to do ever. #ImWithHer"
trvl_god|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
trvl_god|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
stephmarieee|ODOGGOD|0.0|0.0|1.0|0.0|@ODOGGOD same haven't seen one Hillary sign at all
Jessica48911162|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
dallaselaineee|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
lonelyabstract|chasemylovex|-0.3586|0.127|0.873|0.0|"RT @chasemylovex: no, Hillary is not the ""ideal candidate"" but we still gonna vote for her tho... and we'll deal with sis later, ya hear me"
jaqueoozi|ThatKarnMcCloud|0.0|0.0|1.0|0.0|"@ThatKarnMcCloud PAHAHAHA NEVER HEARD THAT GEM OF POLITICAL COMMENTARY BEFORE! HEY KARN, TRUMP HAS GOOFY HAIR AND HILLARY DABBED ONCE! PFFFT"
TuNaLdO|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
TuNaLdO|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
spacesoons|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
knlaguerre|thetrudz|0.0|0.0|1.0|0.0|"RT @thetrudz: History, Symbolism &amp; Representation: Examining The Meaning of Hillary Rodham Clinton's Rise https://t.co/9EPPKpGgKe https://t"
knlaguerre|thetrudz|0.0|0.0|1.0|0.0|"RT @thetrudz: History, Symbolism &amp; Representation: Examining The Meaning of Hillary Rodham Clinton's Rise https://t.co/9EPPKpGgKe https://t"
rodawyd|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
JayMcIntyre1|BobMacAZ|0.2023|0.0|0.904|0.096|"RT @BobMacAZ: CIA Officially Breaks Their Silence, Reveals Top Secret Info on Hillary Shes Done https://t.co/oFQmT2ksXI via @USADailyInfo"
JayMcIntyre1|dailyinfo|0.2023|0.0|0.904|0.096|"RT @BobMacAZ: CIA Officially Breaks Their Silence, Reveals Top Secret Info on Hillary Shes Done https://t.co/oFQmT2ksXI via @USADailyInfo"
JDOZIER66|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
JDOZIER66|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
Jzumble|ReVamPT_EvL|0.0|0.0|1.0|0.0|RT @ReVamPT_EvL: Kids nationwide once Hillary gets in office. Don't let this happen https://t.co/FYJ3I0qaUB
Jzumble|twitter|0.0|0.0|1.0|0.0|RT @ReVamPT_EvL: Kids nationwide once Hillary gets in office. Don't let this happen https://t.co/FYJ3I0qaUB
ajvandenburgh|ConstanceQueen8|0.0|0.0|1.0|0.0|RT @ConstanceQueen8: Tracking Voter TurnOutHope This TrendsIn The Other 44 States#Vote4Trump #Defeat_Hillary#HillaryForPrisi
RyanQC1|LarsLarsonShow|0.0|0.0|1.0|0.0|@LarsLarsonShow driving up to 05 and out patent just now 200 Trump signs not one Hillary
CarolCcsee|MaryLoveUS4|0.4939|0.0|0.833|0.167|RT @MaryLoveUS4: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/br0QOB4q2R https://t
CarolCcsee|thegatewaypundit|0.4939|0.0|0.833|0.167|RT @MaryLoveUS4: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/br0QOB4q2R https://t
ELZUNIA79|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
teameray|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
teameray|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
CalebBrankle|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
CalebBrankle|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
wmhjames|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
wmhjames|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
deryloconstruct|Pamela_Moore13|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
deryloconstruct|twitter|-0.7959|0.415|0.585|0.0|RT @Pamela_Moore13: Indiana is joining Kentucky saying Hell No to Hillary! https://t.co/Ip6DZVgiaa
whomadewho102|HaskelBiz|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
whomadewho102|twitter|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
MiTreasurHunter|twitter|-0.8034|0.341|0.573|0.086|DEMOCRATS are VIOLENT! Got verbally assaulted by a foul mouthed female Hillary supporter today. HILLARY will furthe https://t.co/kLWgh4pY1s
JohnCricket7|perezhilton|0.0|0.0|1.0|0.0|Alec Baldwin And Kate McKinnon Break Character To Knock Some Sense Into America  W https://t.co/x2Y209V2hT
Aubrey_Mays97|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
Aubrey_Mays97|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
cocoapencil101|Lexual__|0.3182|0.0|0.905|0.095|RT @Lexual__: Another comment: all the things y'all mentioned Hillary doing I'm sure Trump would have done if he had a career in politics.
hrh_orchid|robynkanner|0.2103|0.0|0.923|0.077|RT @robynkanner: ***** FLORIDA &amp; NORTH CAROLINA ******POLLS CLOSE SOON. STAY IN LINE. YOUR VOTE FOR HILLARY CLINTON MATTERS SO SO SO SO M
nayteer|summerpennell|0.0|0.0|1.0|0.0|RT @summerpennell: Voting for Hillary with my fellow @UNCAlumni @UNCSchoolofEd professors #ProfessorsInPantsuits #PantsuitNation #We'reWith
petalnh|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
cisppetta|Scarlett210|-0.6597|0.234|0.766|0.0|RT @Scarlett210: If U can vote 4 #Hillary when you KNOW she's seriously ill maybe U shld forget ur enormous #Obamacare payt &amp; go to the hos
AAlanyaodom1|LifeAsRednecks|0.6124|0.0|0.773|0.227|RT @LifeAsRednecks: Votin for Hillary just because shes a woman is like drinkin antifreeze just because it looks like Gatorade.
SON_DJunior|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
BeaThePort|keiradanvers|0.8225|0.0|0.714|0.286|"@keiradanvers @7_MotorSport as they said trump was expected to win those, but hillary will win the big states with most votes"
savyyysav|KayzoMusic|0.765|0.0|0.68|0.32|RT @KayzoMusic: If Hillary Clinton wins I hope she comes out for her victory speech to jotaro.
CRETE288|nytimes|0.2991|0.162|0.577|0.262|@nytimes for sure Hillary Clinton  isn't telling the truth!!!
spookyhan1975|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
SuzieQt154320|1stAirDel_USMCR|-0.1406|0.075|0.925|0.0|"RT @1stAirDel_USMCR: Single mom faces charges for selling home-cooked meals in a Facebook group, but  Hillarys crimes not big enough https"
DonaldB34044603|coachVMarino|0.4404|0.0|0.884|0.116|@coachVMarino @seanhannity I have worked up and down the coast of florida working on boats and nobody had anything good to say about Hillary
spreadthemesg|guntrust|0.0|0.0|1.0|0.0|"RT @guntrust: WikiLeaks:Hillary's campaign wants ""unaware"" and ""compliant"" citizens https://t.co/yRva216Xm4 #tcot #2A #Trump via @guntrust"
spreadthemesg|lawnews|0.0|0.0|1.0|0.0|"RT @guntrust: WikiLeaks:Hillary's campaign wants ""unaware"" and ""compliant"" citizens https://t.co/yRva216Xm4 #tcot #2A #Trump via @guntrust"
CallMeZaaddyyy|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
CallMeZaaddyyy|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
AnnJone70245663|GrrrGraphics|0.0|0.0|1.0|0.0|RT @GrrrGraphics: Ooops! see what @Reuters did! https://t.co/ptfuUrekjX
AnnJone70245663|thegatewaypundit|0.0|0.0|1.0|0.0|RT @GrrrGraphics: Ooops! see what @Reuters did! https://t.co/ptfuUrekjX
taylorsinsanity|agentscullly|-0.2401|0.213|0.633|0.154|RT @agentscullly: I'm not American but honestly scared for u all+the result will have an impact on the whole world so I better wake up to H
apeaceofcake_10|WTF_Eh|0.8442|0.058|0.576|0.366|"RT @WTF_Eh: People tweeting ""pray Hillary wins""  The party that boo's God &amp; removed Him from their platform. Shake my head. #ElectionNight"
lunchbox1034|RealVinnieJames|0.4574|0.0|0.728|0.272|"RT @RealVinnieJames: #WTFAmericaIn5Words - ""Hillary voters support THESE THINGS?!"" https://t.co/NMrdKLJvpX"
lunchbox1034|twitter|0.4574|0.0|0.728|0.272|"RT @RealVinnieJames: #WTFAmericaIn5Words - ""Hillary voters support THESE THINGS?!"" https://t.co/NMrdKLJvpX"
Kashii_Nap|blvckpapii|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
Kashii_Nap|twitter|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
RinsseuxQC|iHateAntony|0.8126|0.0|0.575|0.425|RT @iHateAntony: My face when Trump wins vs when Hillary wins. https://t.co/y2H2XX9LC8
RinsseuxQC|twitter|0.8126|0.0|0.575|0.425|RT @iHateAntony: My face when Trump wins vs when Hillary wins. https://t.co/y2H2XX9LC8
TeddyScibelli|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Barbara40940975|CrappyMovies|-0.296|0.128|0.872|0.0|"RT @CrappyMovies: @realDonaldTrump @CNN oh, in 2004 no one bitched...i got my Hillary vote in https://t.co/ZpUxkCUEcW"
Barbara40940975|twitter|-0.296|0.128|0.872|0.0|"RT @CrappyMovies: @realDonaldTrump @CNN oh, in 2004 no one bitched...i got my Hillary vote in https://t.co/ZpUxkCUEcW"
brianabutcher|BuzzFeed|0.4019|0.0|0.838|0.162|RT @BuzzFeed: People are wearing pantsuits today to show their support for Clinton https://t.co/Tr03g8tcMZ https://t.co/Zdg04j2uhP
brianabutcher|buzzfeed|0.4019|0.0|0.838|0.162|RT @BuzzFeed: People are wearing pantsuits today to show their support for Clinton https://t.co/Tr03g8tcMZ https://t.co/Zdg04j2uhP
ClarissaSchreed|TheDailyShow|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
ClarissaSchreed|cc|0.0|0.0|1.0|0.0|RT @TheDailyShow: Beyonc performs at a Hillary Clinton rally. https://t.co/TCkTVdEWwB https://t.co/Uo18unNpjY
gladiz_h|gaybubs|0.5319|0.0|0.636|0.364|RT @gaybubs: @Calum5SOS YES VOTE FOR HILLARY
holyvanderjesus|kt_taylor17|0.3612|0.0|0.898|0.102|"RT @kt_taylor17: when i wake up in the morning, im praying thata) hillary will be president b) there'll be a steaming plate of katsu next"
bpweise|AGuyNamedNam|0.0|0.0|1.0|0.0|RT @AGuyNamedNam: you know whites and asians can also vote for hillary right rudy https://t.co/Nhi0I7lp6t
bpweise|twitter|0.0|0.0|1.0|0.0|RT @AGuyNamedNam: you know whites and asians can also vote for hillary right rudy https://t.co/Nhi0I7lp6t
jzertuche15|kayleighguad|0.0|0.0|1.0|0.0|@kayleighguad @ShannonPatter34 *Hillary
deadtrbI|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Heathah_|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
lynsicle|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
mati_romaniello|KaivanShroff|0.6705|0.12|0.602|0.278|RT @KaivanShroff: STAY IN LINE until you get to exercise your right to vote. After a year of hatred let's make sure Hillary wins and wins b
MaryRachBailey|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
MaryRachBailey|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
melofidias|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
jl_shepherd|freckledbutt|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
jl_shepherd|twitter|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
bgspalding|Always_Trump|0.3612|0.0|0.878|0.122|RT @Always_Trump: REMINDER: Hillary passes out and gets chucked into a van like a side of beef #HillarysHealth #ElectionDay #Voted #myvote2
tbarksdl|billmaher|-0.8753|0.382|0.574|0.044|"RT @billmaher: Pls vote for Hillary today. Even if you don't like her, its necessary to block a dangerous lunatic ultimate power. #ThisTime"
defminseok|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
arejaayy_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
arejaayy_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
igor_outeiro|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
MeliNicole_xoxo|BJCalvillo|0.0459|0.145|0.737|0.119|RT @BJCalvillo: If I were to vote it would be for Hillary simply because if Trump wins there will be riots and I don't want someone to stea
smitaprakash|BDUTT|0.3182|0.0|0.796|0.204|@BDUTT I'm at Trump zone. I was at Hillary's y'day :-)
RobertKellaghan|FintanCox|0.6597|0.0|0.779|0.221|"RT @FintanCox: Looking at Those exit polls,Hillary looks like she's going to blow trump out,nutty right wing GOP primary voters effectively"
soph2124|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
memereto4|JaredWyand|0.8941|0.0|0.561|0.439|RT @JaredWyand: ALERT: Everyone make sure your vote is placed accurately. Amazing how all these reports favor Hillary.#ElectionDay #Vote
dejean76|Rach_IC|0.4939|0.0|0.833|0.167|RT @Rach_IC: Ugh... More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/R0yTMEIzBb
dejean76|thegatewaypundit|0.4939|0.0|0.833|0.167|RT @Rach_IC: Ugh... More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/R0yTMEIzBb
LyndaKelly|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
LyndaKelly|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
miladysdewinter|DanaSchwartzzz|0.6249|0.075|0.712|0.214|RT @DanaSchwartzzz: Dear lord if Hillary Clinton wins I'll read a book before bed and stop tweeting so much and give more to the homeless a
AllieGoertz|twitter|-0.5574|0.545|0.455|0.0|Nasty for Hillary  https://t.co/nUrnSjDvDY
higginskiara|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
higginskiara|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
passcon93|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
passcon93|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
MDaviot|lgmaterna|-0.4939|0.132|0.868|0.0|"RT @lgmaterna: #ImVotingBecause Hillary has bombed more children than she has helped, and Bill has jailed more black Americans than he has"
xPLOCC|AthenaElias|0.0|0.0|1.0|0.0|@AthenaElias @DrPresidentPat @realDonaldTrump @EricTrump and Hillary wouldn't ?
mrred549|Pamela_Moore13|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
mrred549|twitter|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
yurbaink|cnni|0.6369|0.0|0.833|0.167|"RT @cnni: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/0RU6ozSJGg"
yurbaink|cnn|0.6369|0.0|0.833|0.167|"RT @cnni: Married for 37 years. He's voting for Hillary. She's voting for Trump. But in the end, there's still love https://t.co/0RU6ozSJGg"
omar_anwari|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
choosycharles|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
choosycharles|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
keycieraa|PETTYMAMII|-0.8441|0.269|0.731|0.0|RT @PETTYMAMII: Vote Hillary Clinton idc is she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
IrcinkSuzanne|KingAJ40|0.6209|0.0|0.747|0.253|RT @KingAJ40: Good People of MICHIGAN!!! Don't Let Hillary Clinton CONFISCATE your GUNS!!!https://t.co/E7zbgg966nhttps://t.co/I97WEXYJNE
IrcinkSuzanne|t|0.6209|0.0|0.747|0.253|RT @KingAJ40: Good People of MICHIGAN!!! Don't Let Hillary Clinton CONFISCATE your GUNS!!!https://t.co/E7zbgg966nhttps://t.co/I97WEXYJNE
RileyKaftonn|twitter|0.0|0.0|1.0|0.0|When someone says they're voting for Hillary https://t.co/Ynu9eY6mpB
BabyMattss|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
BabyMattss|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
sophieissoapy|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
sophieissoapy|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
ramirezlisully|NasMaraj|0.0|0.0|1.0|0.0|"RT @NasMaraj: If this doesn't make you vote Hillary, I don't know what will. #ImWithHer https://t.co/shQYaBFeGR"
ramirezlisully|twitter|0.0|0.0|1.0|0.0|"RT @NasMaraj: If this doesn't make you vote Hillary, I don't know what will. #ImWithHer https://t.co/shQYaBFeGR"
nohelyshoot|cammiescott|0.3612|0.0|0.783|0.217|RT @cammiescott: Like for Hillary. Retweet for Hillary.(unfollow for Trump)
tarahgeeface|Lanniyahh|0.5719|0.0|0.764|0.236|RT @Lanniyahh: &amp;I I'm wearing my sticker to work tmrw when Hillary wins 
Harneil_A|twitter|0.3818|0.1|0.704|0.196|... a media outlet that is in favour of trump could make a list for Hillary too. Media fooling people too easily th https://t.co/QKBpzGy0Kz
leonela_xo|meechonmars|0.3612|0.0|0.909|0.091|RT @meechonmars: voting for hillary when you wanted to vote for bernie is like when you ask for a coke and they say they have pepsi products
J_JonesIV|michaelharrisII|-0.5106|0.155|0.845|0.0|RT @michaelharrisII: The thought of Hillary Clinton being elected president tomorrow night literally makes me sick to my stomach
badgalkekeee|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
badgalkekeee|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
lizthemermaid|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
lizthemermaid||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
Worped4|HAGOODMANAUTHOR|0.9474|0.0|0.525|0.475|RT @HAGOODMANAUTHOR: TRUMP WINS FLORIDA!!! TRUMP WINS FLORIDA!!! TRUMP WINS FLORIDA!! (Remember when they'd call a state for Hillary over B
stevuhn1027|austinn_holland|-0.5291|0.424|0.576|0.0|RT @austinn_holland: Hillary sucks but not like Monica
tay_rizzuto|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
tay_rizzuto|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
FewerHorsesNBay|MakeupArtistmag|0.0|0.0|1.0|0.0|RT @MakeupArtistmag: We're voting for the 'SNL' make-up/hair team for their Hillary Clinton and Donald Trump transformations! https://t.co/
FewerHorsesNBay|t|0.0|0.0|1.0|0.0|RT @MakeupArtistmag: We're voting for the 'SNL' make-up/hair team for their Hillary Clinton and Donald Trump transformations! https://t.co/
styinyoureye|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
styinyoureye|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
fuckoffbeth|yvezayntIaurent|-0.5423|0.22|0.78|0.0|"RT @yvezayntIaurent: white person: idk whos worse: hillary or trumplgbtq, women, black people, immigrants, muslims: trump iswhite pers"
Nellie20K|michaelbeatty3|0.0|0.0|1.0|0.0|RT @michaelbeatty3: GOLDMAN SACHS SCRIPTED ANSWERS?#Hillary #FeelTheBern #CNN  #PodestaEmails35 #Wikileaks #electionday https://t.co/
Nellie20K|t|0.0|0.0|1.0|0.0|RT @michaelbeatty3: GOLDMAN SACHS SCRIPTED ANSWERS?#Hillary #FeelTheBern #CNN  #PodestaEmails35 #Wikileaks #electionday https://t.co/
Goodnightma|LastWave2014|-0.3818|0.191|0.809|0.0|"RT @LastWave2014: Media lied, Bush DID NOTE vote for Hillary Clinton https://t.co/SWf3EmjXyz"
Goodnightma|nbcconnecticut|-0.3818|0.191|0.809|0.0|"RT @LastWave2014: Media lied, Bush DID NOTE vote for Hillary Clinton https://t.co/SWf3EmjXyz"
ashhley33|JLaughmiller|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
ashhley33|twitter|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
Reesesuth|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
tinaapratt|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
Jeancarlos_GC|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
blackle0patra|Lexual__|0.3182|0.0|0.905|0.095|RT @Lexual__: Another comment: all the things y'all mentioned Hillary doing I'm sure Trump would have done if he had a career in politics.
Kardorian79|mitchellvii|-0.3182|0.206|0.653|0.141|"RT @mitchellvii: If true, this is brutal for Hillary.  She won't match Obama's numbers. https://t.co/z0o069Bv1p"
Kardorian79|twitter|-0.3182|0.206|0.653|0.141|"RT @mitchellvii: If true, this is brutal for Hillary.  She won't match Obama's numbers. https://t.co/z0o069Bv1p"
bradymyers32|ChaseMatthews98|0.5267|0.0|0.764|0.236|RT @ChaseMatthews98: Hillary's winning because all of the republicans are out working
BordersAreGreat|HuffingtonPost|-0.34|0.124|0.876|0.0|@HuffingtonPost has shamelessly campaigned for corrupt Hillary. 1st time in 20 years we've had possibility of REAL https://t.co/ISQcGfbX0i
BordersAreGreat|twitter|-0.34|0.124|0.876|0.0|@HuffingtonPost has shamelessly campaigned for corrupt Hillary. 1st time in 20 years we've had possibility of REAL https://t.co/ISQcGfbX0i
GeorgiaDaskalos|DRUDGE_REPORT|0.3182|0.0|0.827|0.173|RT @DRUDGE_REPORT: Madonna breaks promise to give oral to Hillary voters... https://t.co/obsQ3RlTFO
GeorgiaDaskalos|nydailynews|0.3182|0.0|0.827|0.173|RT @DRUDGE_REPORT: Madonna breaks promise to give oral to Hillary voters... https://t.co/obsQ3RlTFO
DelawareFreedom|newsmax|0.4404|0.0|0.734|0.266|RT @newsmax: Unpredictable Trump Better Than Scandal-laden Hillary  https://t.co/8DABeBwZVo
DelawareFreedom|newsmax|0.4404|0.0|0.734|0.266|RT @newsmax: Unpredictable Trump Better Than Scandal-laden Hillary  https://t.co/8DABeBwZVo
SandyCharara|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
SandyCharara|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
sadgallexi|twitter|-0.5106|0.155|0.845|0.0|"""Hillary is a liar, listen to me while I parrot things people have been saying for years to sound smart."" https://t.co/sN2AxnIpbD"
good4politics|jmartNYT|0.0|0.0|1.0|0.0|@jmartNYT @R_Love317 I saw other tweets claiming they voted for Hillary
TheNikkiG|emerylord|0.2023|0.09|0.789|0.12|RT @emerylord: listen I know she's not Obama in terms of firing people up...but Hillary inspired a bunch of WRITERS to put on PANTS today..
spain_zoe|diiegooo94|0.0|0.0|1.0|0.0|"RT @diiegooo94: If Hillary gets Elected I'm not coming to school, if they file truancy on me I will state""If our president can break the la"
KaineMilner_|HillaryClinton|0.0|0.0|1.0|0.0|Come on Hillary!! #FuckTrump #ImWithHer @HillaryClinton
a4beach|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
SalmaBar|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
SalmaBar|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
JaredStrackbein|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
BarbaraZaccai|mitchellvii|-0.7003|0.225|0.775|0.0|"RT @mitchellvii: Based upon what I am seeing from Tampa and numbers have remained stead all day, Hillary will lose Florida and badly."
tomasnjill|CalmNcanny|0.7199|0.0|0.807|0.193|@CalmNcanny NOPE! AND I WENT THERE TWICE THIS YEAR TO EDUCATE THEM AND THEY AREN'T VOTING ! THEY OWN HILLARY'S POLICY IF SHE WINS.
DarriusKV|twitter|0.0772|0.0|0.86|0.14|"Vote for who you want, vote for Hillary https://t.co/oxGyhowtEt"
h_blundell|twitter|0.4404|0.0|0.879|0.121|I hope I am going to wake up and see millions of tweets about Hillary Clinton being the next President or my expres https://t.co/evkL6fVMB2
AyawnuhMayree|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
AyawnuhMayree|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Mangoluu|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
sebastianchiap|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
OccuWorld|infiniteunknown|0.0|0.0|1.0|0.0|68% Of Saudis Prefer Hillary Clinton As U.S. President https://t.co/d2OL6GHPR8
GFabrygherardi|GMA|0.0|0.0|1.0|0.0|"RT @GMA: ""All Hillary Clinton needs to do is hold all of the states where she currently has a lead."" - @jonkarl https://t.co/OwlrhGvIKj"
GFabrygherardi|twitter|0.0|0.0|1.0|0.0|"RT @GMA: ""All Hillary Clinton needs to do is hold all of the states where she currently has a lead."" - @jonkarl https://t.co/OwlrhGvIKj"
gkoogz|ConstanceQueen8|0.0|0.0|1.0|0.0|RT @ConstanceQueen8: Tracking Voter TurnOutHope This TrendsIn The Other 44 States#Vote4Trump #Defeat_Hillary#HillaryForPrisi
honradojhuztin|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
jrbixby|PrisonPlanet|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
jrbixby|pittsburgh|0.4404|0.0|0.838|0.162|RT @PrisonPlanet: Trump supporters in Pennsylvania seeing their votes switched to Hillary before their eyes. https://t.co/hfgye7AKaJ
changeisneeded_|BlissTabitha|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
changeisneeded_|weaselzippers|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
Navyboy08021|AbbyMartinM|-0.3182|0.228|0.642|0.13|"RT @AbbyMartinM: Colin Powell TRUTH Revealed In Last Moments, Hillary Used Obama To HIDE Her Treason https://t.co/WutfwCHhkg https://t.co/E"
Navyboy08021|endingthefed|-0.3182|0.228|0.642|0.13|"RT @AbbyMartinM: Colin Powell TRUTH Revealed In Last Moments, Hillary Used Obama To HIDE Her Treason https://t.co/WutfwCHhkg https://t.co/E"
Jamesmel|DVATW|0.5106|0.0|0.87|0.13|RT @DVATW: Bill Clinton tried to cheer up Hillary today by reminding her that Mandela wasn't elected president until after serving 27 yrs i
superdryhowell|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
superdryhowell|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
haleeshiann|AllisonRenee_14|0.7391|0.0|0.734|0.266|RT @AllisonRenee_14: Collin was born @ 35wks and is perfectly healthy but Hillary Clinton thinks its ok to have abortions all the way till
_bayelizabeth_|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
BrextonIsaacs|kylegriffin1|0.6369|0.0|0.846|0.154|"RT @kylegriffin1: Clinton camp out w/ new behind-the-scenes vids of HRC, best may be Bill jumping up and down after the 1st debate: https:/"
BrextonIsaacs||0.6369|0.0|0.846|0.154|"RT @kylegriffin1: Clinton camp out w/ new behind-the-scenes vids of HRC, best may be Bill jumping up and down after the 1st debate: https:/"
ChrisGiamatti|umpire43|0.0|0.0|1.0|0.0|RT @umpire43: A woman in Fla reported she voted Trump on Smartmatic https://t.co/Sm6mmsb0AH was flipped to Hillary and multiplied to 200 in
ChrisGiamatti||0.0|0.0|1.0|0.0|RT @umpire43: A woman in Fla reported she voted Trump on Smartmatic https://t.co/Sm6mmsb0AH was flipped to Hillary and multiplied to 200 in
Hideyoshi_Lover|wendeezyv2|-0.8402|0.45|0.55|0.0|@wendeezyv2 @fuckinweeb hillary is sakura becauses she is ugly useless and everybody hates her
M_i_r_e_y_a_|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
M_i_r_e_y_a_|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
sandra79707|Scarlett210|-0.6597|0.234|0.766|0.0|RT @Scarlett210: If U can vote 4 #Hillary when you KNOW she's seriously ill maybe U shld forget ur enormous #Obamacare payt &amp; go to the hos
BestWebEnglish|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
BestWebEnglish|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
nitroman05|bry_shook|-0.5106|0.231|0.769|0.0|@bry_shook @HillaryClinton  the whole thing is a joke.. hillary should be in prison
goghstly|PoeticsNormani|0.7717|0.0|0.309|0.691|RT @PoeticsNormani: Hillary better win
suidfc|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/FbSc1sQ8jN
suidfc|nbcconnecticut|0.0|0.0|1.0|0.0|I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news. https://t.co/FbSc1sQ8jN
MatthewMcM23|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
MatthewMcM23|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
soccer_sara13|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
soccer_sara13|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
josephiykech|sheila06942158|-0.3382|0.123|0.877|0.0|"RT @sheila06942158: While Polls are Still Open, FBI Agents Drop the Biggest Bombshell Ever on HILLARY CLINTON! https://t.co/anDXtdOsSR"
josephiykech|lsh|-0.3382|0.123|0.877|0.0|"RT @sheila06942158: While Polls are Still Open, FBI Agents Drop the Biggest Bombshell Ever on HILLARY CLINTON! https://t.co/anDXtdOsSR"
DemencjuszX|Daily_Express|-0.2263|0.159|0.725|0.116|RT @Daily_Express: Voter's angry response after being asked if she was excited about Clinton becomming president #USElection2016https://t.
BethHawkins10|BruceBartlett|0.6311|0.076|0.688|0.235|"RT @BruceBartlett: For the record, I voted enthusiastically for Hillary Clinton today. She may not be perfect, but she's light years better"
dtav|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
dtav|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
cessjet|HaskelBiz|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
cessjet|twitter|0.128|0.127|0.724|0.149|RT @HaskelBiz: India Smith voted for Trump because Hillary Clinton 'broke the trust of the country' #haelex https://t.co/J0LAqXacli
oneideatoday|giphy|0.5859|0.0|0.787|0.213|"New trending GIF tagged loop, donald trump, hillary clinton, winner, trump v clinton via G https://t.co/T6nKKblVd7 https://t.co/ur5FX9u5mf"
slkn11|geoffgarin|0.5423|0.0|0.816|0.184|"RT @geoffgarin: I am going to be ecstatic when Hillary Clinton wins tonight.  Not just because Trump won't be president, but more because s"
HunterC_3|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
Quack4Bernie|wikileaks|-0.2732|0.139|0.861|0.0|RT @wikileaks: Its ignorant to vote for Hillary Clinton without reading WikiLeaks https://t.co/Tiywc9Nrgr https://t.co/c0QaJW4hCi
Quack4Bernie|denverpost|-0.2732|0.139|0.861|0.0|RT @wikileaks: Its ignorant to vote for Hillary Clinton without reading WikiLeaks https://t.co/Tiywc9Nrgr https://t.co/c0QaJW4hCi
meghanxokate|nationdivided|-0.68|0.248|0.665|0.087|"RT @nationdivided: Very first results is in, thank you Kentucky Coal Country says Hell no to Hillary! Go Trump #MAGS #Election2016 https://"
meghanxokate||-0.68|0.248|0.665|0.087|"RT @nationdivided: Very first results is in, thank you Kentucky Coal Country says Hell no to Hillary! Go Trump #MAGS #Election2016 https://"
vincentcasanov1|fuckinfenty|-0.5719|0.252|0.748|0.0|RT @fuckinfenty: Me: I hate Hillary Clinton Rihanna: wears Hillary Clinton shirtMe: https://t.co/bkUXzFP68Z
vincentcasanov1|twitter|-0.5719|0.252|0.748|0.0|RT @fuckinfenty: Me: I hate Hillary Clinton Rihanna: wears Hillary Clinton shirtMe: https://t.co/bkUXzFP68Z
crime18458238|WordSmithGuy|0.7595|0.0|0.705|0.295|"RT @WordSmithGuy: Pennsylvania, Ohio &amp; Michigan Voters: Remember how little Hillary cares about the Clean Coal Industry. VOTE for Energy In"
kathewineposada|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
kathewineposada|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
SuzannaChaparro|cursedsalad|-0.1007|0.18|0.663|0.157|RT @cursedsalad: Electoral College is refusing to accept Hillary's corruption! #RestoreChecksandBalances #ElectionNight #WTFAmericaIn5Words
derrickraju66|IngrahamAngle|0.0|0.0|1.0|0.0|RT @IngrahamAngle: Hillary needs celebs to draw crowds. Trump doesn't. He has an actual plan to grow jobs &amp; enforce rule of law. https://t.
derrickraju66||0.0|0.0|1.0|0.0|RT @IngrahamAngle: Hillary needs celebs to draw crowds. Trump doesn't. He has an actual plan to grow jobs &amp; enforce rule of law. https://t.
ThomasCayo1|WeNeedTrump|0.0|0.0|1.0|0.0|RT @WeNeedTrump: Twitter wants Donald Trump. 264K retweets for Donald Trump. 35.6K retweets for Hillary Clinton. #MakeAmericaGreatAgain htt
maryjanerdz1103|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
maryjanerdz1103|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Wambamphilosoph|KrackKids|0.0|0.0|1.0|0.0|RT @KrackKids:  When you have to vote for Trump or Hillary. https://t.co/VJyfkSbTKp
Wambamphilosoph|vine|0.0|0.0|1.0|0.0|RT @KrackKids:  When you have to vote for Trump or Hillary. https://t.co/VJyfkSbTKp
laura_paredess|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
LackneyMichelle|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
LackneyMichelle|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
tsuttonNYC|billmaher|-0.8753|0.382|0.574|0.044|"RT @billmaher: Pls vote for Hillary today. Even if you don't like her, its necessary to block a dangerous lunatic ultimate power. #ThisTime"
lashingsoflove|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
lashingsoflove|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
shershul_|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
shershul_|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
t_moneeeyyyy|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
t_moneeeyyyy|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
RickTheGeneral|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
RickTheGeneral|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
ChuckNoyes|AbbyMartin|-0.6423|0.258|0.645|0.097|@AbbyMartin  Libya did not attack us . 90% of casualties in Modern War are WOMEN  and children..who hates women mor https://t.co/zuHsDnDbqa
ChuckNoyes|twitter|-0.6423|0.258|0.645|0.097|@AbbyMartin  Libya did not attack us . 90% of casualties in Modern War are WOMEN  and children..who hates women mor https://t.co/zuHsDnDbqa
PatriotinMO_USA|LifeZette|0.4404|0.0|0.791|0.209|RT @LifeZette: Why @realDonaldTrump would be a better president for American women https://t.co/dyLBBgeB2c
PatriotinMO_USA|lifezette|0.4404|0.0|0.791|0.209|RT @LifeZette: Why @realDonaldTrump would be a better president for American women https://t.co/dyLBBgeB2c
RealTimeHack|nytimes|0.0|0.0|1.0|0.0|How the FBI Reviewed Thousands of Emails in One Week - New York Times https://t.co/utgnyG6CHu #GN
FeeElleby|NasMaraj|0.0|0.0|1.0|0.0|"RT @NasMaraj: If this doesn't make you vote Hillary, I don't know what will. #ImWithHer https://t.co/shQYaBFeGR"
FeeElleby|twitter|0.0|0.0|1.0|0.0|"RT @NasMaraj: If this doesn't make you vote Hillary, I don't know what will. #ImWithHer https://t.co/shQYaBFeGR"
scottishphoenix|Mrs_KittyO|0.0|0.0|1.0|0.0|@Mrs_KittyO Will I be able to resist being naughty and mischievous tonight on here if Hillary wins?! 
andrewkmorse|CNET|0.0|0.0|1.0|0.0|Can social media call the election? https://t.co/mh9iX9EXCD via @CNET #Election2016 #ElectionNight
andrewkmorse|cnet|0.0|0.0|1.0|0.0|Can social media call the election? https://t.co/mh9iX9EXCD via @CNET #Election2016 #ElectionNight
sheila06942158|TRay1949|0.0|0.0|1.0|0.0|RT @TRay1949: Hillary's Kissin KKK  https://t.co/2RoehKOfht
sheila06942158|twitter|0.0|0.0|1.0|0.0|RT @TRay1949: Hillary's Kissin KKK  https://t.co/2RoehKOfht
_JasonAA|Poochda63|0.3948|0.079|0.777|0.144|RT @Poochda63: Don't play with me I'll show up knocking RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
DougNelson48|YouTube|0.0|0.0|1.0|0.0|"Julian Assange just did it: WikiLeaks Dispenses 23,000 MORE Hillary Em... https://t.co/4joZ2LZPs0 via @YouTube"
DougNelson48|youtube|0.0|0.0|1.0|0.0|"Julian Assange just did it: WikiLeaks Dispenses 23,000 MORE Hillary Em... https://t.co/4joZ2LZPs0 via @YouTube"
cfsuburbia|PopCrave|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
cfsuburbia|twitter|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
bodyblissbyj|kle317|0.0|0.0|1.0|0.0|@kle317 @Brian_Pilgrim40 Bloomberg is in bed with Hillary...not credible
WUTWNG91|_donaldson|0.3182|0.0|0.85|0.15|@_donaldson @rickhasen @joshtpm so these blacks on a church bus is responsible for a Hillary email?
BettyGebruu|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
BettyGebruu|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Oldstones70|Delo_Taylor|0.0|0.0|1.0|0.0|RT @Delo_Taylor: Side note: Hillary Clinton is White. https://t.co/J0QdqGRv5v
Oldstones70|twitter|0.0|0.0|1.0|0.0|RT @Delo_Taylor: Side note: Hillary Clinton is White. https://t.co/J0QdqGRv5v
Shalom555222|mitchellvii|-0.7645|0.32|0.68|0.0|"RT @mitchellvii: Based upon exits, voters very unhappy with big money corruption.  That's bad for Hillary."
Baddicey|twitter|-0.347|0.213|0.787|0.0|Anywho... DO IT FA HILLARY SHAKE IT FA HILLARY https://t.co/yg5V2PATle
venzuelanprince|Madonna|0.8877|0.0|0.605|0.395|RT @Madonna: Last night was. Amazing!!! Save this Country please!!  Vote for Hillary Clinton!  Today is the Day!  https://t
venzuelanprince||0.8877|0.0|0.605|0.395|RT @Madonna: Last night was. Amazing!!! Save this Country please!!  Vote for Hillary Clinton!  Today is the Day!  https://t
RolandoMederos|FoxNews|0.3182|0.0|0.777|0.223|@FoxNews @realDonaldTrump @HillaryClinton fuc.... Hillary. .please lord go Trump
CALIFUK|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
roykolepoyko|markhumphrys|-0.2023|0.079|0.921|0.0|"@markhumphrys in fact, trump is closer to marxism than hillary. left &amp; right people are often unaware fascism started from national plebeian"
arierango|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
lifeliner2|billmaher|-0.8753|0.382|0.574|0.044|"RT @billmaher: Pls vote for Hillary today. Even if you don't like her, its necessary to block a dangerous lunatic ultimate power. #ThisTime"
shirleycolleen|BlissTabitha|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
shirleycolleen|weaselzippers|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
blooprr|WikiLeaksParty|0.0|0.0|1.0|0.0|@WikiLeaksParty Especially when Hillary takes over. Podesta's mouth will be watering #CheesPizza
jmatz10|WTF_Eh|0.8442|0.058|0.576|0.366|"RT @WTF_Eh: People tweeting ""pray Hillary wins""  The party that boo's God &amp; removed Him from their platform. Shake my head. #ElectionNight"
sanhasflowers|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
HANN_itToAh|chungaah|0.3818|0.122|0.667|0.211|RT @chungaah: Not even worried about the election Ik who gonna win Hillary obviously 
bneil_3|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
bneil_3|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
Antbob_Drums|Liberienne|0.34|0.112|0.68|0.208|RT @Liberienne: Y'all ready for Bill Clinton to be the first lady? Hopefully Hillary cheats on him while in office.
MasonDeVries5|brennan_moody3|0.5719|0.0|0.748|0.252|RT @brennan_moody3: This country will take the fattest L if Hillary wins tonight.
starboyissa|twitter|0.0|0.0|1.0|0.0|why did I get Hillary https://t.co/M0wch2nxgj
esonino|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Jshen2014365|RobWolf_|0.0772|0.0|0.947|0.053|"@RobWolf_ @Bookieinsiders can't see Hillary not taking Florida, Latinos out in big number similar to blacks in 08 and we know what that mean"
kincannon_show|SLandinSoCal|0.0|0.0|1.0|0.0|RT @SLandinSoCal: Does #Hillary have #Kuru? Contracted through #Canabalism. Symptoms mimic #Parkinsons. Would explain her inappropriate out
dejaharianna|thecityofjules|0.4767|0.106|0.683|0.212|RT @thecityofjules: me preparing my fake smile for when hillary wins and white women start talkin bout how far the suffragettes have come h
EastVillageYYC|twitter|-0.2235|0.09|0.91|0.0|Repost from #OutsidersRunClub. Hillary and Trump are in the running tonight - why not join 'em? Run starts at 6:30p https://t.co/SRSARb4jG3
nadiaissocool|vickto_willy|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
nadiaissocool|t|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
_LookDontTouch|Empress_Orit|0.7184|0.216|0.448|0.336|"RT @Empress_Orit: There's BLACK Women stomping hard for Hillary but refused to support or amplify any legit BLACK freedom fighter, fighting"
Urbann_Flora|NasMaraj|0.0|0.0|1.0|0.0|"RT @NasMaraj: If this doesn't make you vote Hillary, I don't know what will. #ImWithHer https://t.co/shQYaBFeGR"
Urbann_Flora|twitter|0.0|0.0|1.0|0.0|"RT @NasMaraj: If this doesn't make you vote Hillary, I don't know what will. #ImWithHer https://t.co/shQYaBFeGR"
presswiz|TheEconomist|0.0762|0.0|0.933|0.067|RT @TheEconomist: The next president will be either Donald Trump or Hillary Clinton. The choice is not hard https://t.co/bInZYYXeW8
presswiz|twitter|0.0762|0.0|0.933|0.067|RT @TheEconomist: The next president will be either Donald Trump or Hillary Clinton. The choice is not hard https://t.co/bInZYYXeW8
bonniebethdail3|ConstanceQueen8|0.0|0.0|1.0|0.0|RT @ConstanceQueen8: Tracking Voter TurnOutHope This TrendsIn The Other 44 States#Vote4Trump #Defeat_Hillary#HillaryForPrisi
nancyl367|worldnetdaily|0.516|0.0|0.836|0.164|"RT @worldnetdaily: CHURCH TAKES BOLD, ANTI-HILLARY STANCEPastor willing to give anyone a ride to polls, irrespective of vote https://t.co"
nancyl367|t|0.516|0.0|0.836|0.164|"RT @worldnetdaily: CHURCH TAKES BOLD, ANTI-HILLARY STANCEPastor willing to give anyone a ride to polls, irrespective of vote https://t.co"
lesdotcomm|michelleelopz|0.5859|0.0|0.798|0.202|RT @michelleelopz: Leslie isn't voting because she saw a tweet that Hillary is going to win  https://t.co/Aj3Fr3zsWC
lesdotcomm|twitter|0.5859|0.0|0.798|0.202|RT @michelleelopz: Leslie isn't voting because she saw a tweet that Hillary is going to win  https://t.co/Aj3Fr3zsWC
mrburlesk|twitter|-0.4767|0.147|0.853|0.0|#FascinatingIf I were Hillary I would be fake ordering bunches of pizzas to be sent to the Trump campaign HQ. https://t.co/sgbF39u3Ns
KGBVeteran|FoxNews|0.7804|0.0|0.605|0.395|@FoxNews is saying that GA and TX are in play for Hillary. This is a joke.
FedoraPayan|RhondaRehbein|0.7579|0.0|0.683|0.317|RT @RhondaRehbein: Pat Buchanan Says The Country Will Not Be United If Hillary Wins | enVolve https://t.co/jXN3fU5wkl
FedoraPayan|en-volve|0.7579|0.0|0.683|0.317|RT @RhondaRehbein: Pat Buchanan Says The Country Will Not Be United If Hillary Wins | enVolve https://t.co/jXN3fU5wkl
_Reagannn|kiingdarry|0.6249|0.102|0.665|0.232|"RT @kiingdarry: all y'all saying y'all not voting b/c y'all don't believe in Hillary nor Trump, if trump wins Y'ALL BETTER NOT COMPLAIN ABO"
Dadah___|AfroGumOfficiaI|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
Dadah___|twitter|0.0|0.0|1.0|0.0|RT @AfroGumOfficiaI: Hillary Clinton doing the #MannequinChallenge on #ElectionDay  https://t.co/fGOnNfYXWQ
schoremis1|Scarlett210|-0.765|0.28|0.72|0.0|"RT @Scarlett210: And #Hillary is a self-serving #elitist who'll continue #globalist policies, destroy ur safety&amp; deprive ur kids of a futur"
Lez_Brarian|twitter|-0.4767|0.162|0.838|0.0|"Yo, Hillary herself left this note in Pantsuit Nation and I'm crying on the subway #ImWithHer https://t.co/nrLtr3tGhB"
ansleyegarland|kaylaaluke|0.8126|0.0|0.575|0.425|RT @kaylaaluke: me when trump wins vs me when hillary wins https://t.co/MoA58nnhfo
ansleyegarland|twitter|0.8126|0.0|0.575|0.425|RT @kaylaaluke: me when trump wins vs me when hillary wins https://t.co/MoA58nnhfo
eddiegrode78|TheWizKhalifa|-0.9022|0.41|0.59|0.0|RT @TheWizKhalifa: People hate Trump because the media made them hate Trump.People hate Hillary because they are paying attention.#Elec
cliff_helton24|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
DannyChallenger|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
TacticalNewsGuy|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
TacticalNewsGuy|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
skylarariannaa|MTVstyle|0.0|0.0|1.0|0.0|RT @MTVstyle: Rihanna wore a t-shirt of HERSELF wearing a Hillary Clinton t-shirt because SHE IS THE STYLE ICON OUR NATION NEEDS:https://
skylarariannaa||0.0|0.0|1.0|0.0|RT @MTVstyle: Rihanna wore a t-shirt of HERSELF wearing a Hillary Clinton t-shirt because SHE IS THE STYLE ICON OUR NATION NEEDS:https://
jooilong|Daily_Expresshttps//t.co/Rx5RvjWPii|0.0|0.0|1.0|0.0|Only pollsters to get Brexit right say its TRUMP for the White House | @Daily_Expresshttps://t.co/Rx5RvjWPii
PhilKnudsen|hickforco|0.4767|0.0|0.86|0.14|@hickforco Just sent a tweet asking me and five of my friends to vote for Hillary and Democrats down the ballot.
ashlleymaries|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
Paperpennn|Orgetorix|0.0|0.0|1.0|0.0|RT @Orgetorix: America decides: Donald Trump or Hillary Clinton https://t.co/cbHeY8gzZn via @smh
Paperpennn|smh|0.0|0.0|1.0|0.0|RT @Orgetorix: America decides: Donald Trump or Hillary Clinton https://t.co/cbHeY8gzZn via @smh
MrPolishedTfUp|jozenc|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
MrPolishedTfUp|twitter|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
thtman_rell|minajsinner|-0.1779|0.086|0.914|0.0|RT @minajsinner: Do it for Hillary Shake it for Hillary Vote for Hillary Do it for the Clintons https://t.co/7MgtCLiigx
thtman_rell|twitter|-0.1779|0.086|0.914|0.0|RT @minajsinner: Do it for Hillary Shake it for Hillary Vote for Hillary Do it for the Clintons https://t.co/7MgtCLiigx
LeeBrocklebank|_actually_ash|-0.6473|0.265|0.592|0.144|RT @_actually_ash: Oh so youre worried about how Trump talks about women but not how Hillary COVERED UP A YOUNG WOMANS RAPE AND LAUGHED ABO
olaftulen|Ekatherene|0.0|0.0|1.0|0.0|"RT @Ekatherene: @mitchellvii @MarianneHaran Las Vegas has Hillary down by 7% , last night she was down 5%...."
_casketpretty|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
devmoeller|HuggiesD|-0.8779|0.502|0.349|0.149|RT @HuggiesD: Man I didn't vote but I sure as hell hope Hillary doesn't win 
smhrache|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
DeejDelRey|aVeryRichBitch_|0.0|0.0|1.0|0.0|RT @aVeryRichBitch_: She out here making people vote for Hillary LMFAOO https://t.co/8PfhJL8cQk
DeejDelRey|twitter|0.0|0.0|1.0|0.0|RT @aVeryRichBitch_: She out here making people vote for Hillary LMFAOO https://t.co/8PfhJL8cQk
ILoveBernie1|twitter|-0.8689|0.353|0.647|0.0|"Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, https://t.co/T3eGu54ype"
jackie_celeste|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
mikey30nv|dforthof|0.4404|0.0|0.674|0.326|@dforthof is that good news for Hillary
emiliana26|Americooligan|0.0|0.0|1.0|0.0|"RT @Americooligan: Trump up 70.5% to Hillary's 25.8% in Indiana. 35,646 votes to 13,049 (1% reporting). #ElectionNight"
ScottItIs|RepCoriFournier|0.0|0.0|1.0|0.0|RT @RepCoriFournier: This is what @CNN is counting on with the BIG push on their network that Republicans will be voting HILLARY n republic
AnimatorsPal|aulty|0.5859|0.0|0.759|0.241|"RT @aulty: #gif #animation loop, donald trump, hillary clinton, winner, trump v clinton https://t.co/yDUv4Ltg0O"
AnimatorsPal|twitter|0.5859|0.0|0.759|0.241|"RT @aulty: #gif #animation loop, donald trump, hillary clinton, winner, trump v clinton https://t.co/yDUv4Ltg0O"
mommatt27|DrMartyFox|-0.296|0.121|0.879|0.0|RT @DrMartyFox: #ImVotingBecause We Must Stop DUAL #JUSTICEWhere #Deplorables Must Follow The #RuleOfLawWhile #Hillary &amp; Her Cronies
NarrendraM||0.0|0.0|1.0|0.0|"#Republicans are leading in the #Congress elections in #Kentucky, #Indiana https://t.co/lzvX1xTPoT https://t.co/v1RD3nFjtd"
RealTimeHack|usatoday|0.197|0.0|0.871|0.129|Hillary Clinton calls voting for herself a 'most humbling feeling' - USA TODAY https://t.co/gV7BfjE8fp #GN
LyndaKelly|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
LyndaKelly|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1% reporting in Indiana: Trump: 69.52%  Hillary 26.78%https://t.co/gEj5j7aP5X #ElectionNight https://t.co/C7hORH
ThomasBialek2|RealVinnieJames|0.0|0.0|1.0|0.0|"RT @RealVinnieJames: TRUMP VOTERS: NOTE! When early counts show Hillary up, they'll  announce the state for her to get you to think all is"
1stTimeVoter216|1stTimeVoter216|0.25|0.0|0.905|0.095|RT @1stTimeVoter216: Crooked Hillary will forever chance the demographic of America by allowing endless amount of illegals &amp; refugees in. V
soIndi|RicheyCollazo|0.8356|0.0|0.603|0.397|RT @RicheyCollazo: white women: Hillary Clintons win is a win for women!me: WHICH WOMEN?  https://t.co/FONDX957Gy
soIndi|twitter|0.8356|0.0|0.603|0.397|RT @RicheyCollazo: white women: Hillary Clintons win is a win for women!me: WHICH WOMEN?  https://t.co/FONDX957Gy
AchmarBinSchibi|suebell49|-0.2023|0.112|0.816|0.071|@suebell49 Hillary admitted in her paid speeches the No Fly Zone would require the deaths of many Syrians
DubWeyer|twitter|-0.5423|0.123|0.877|0.0|When people say they voted for Hillary just BC she is a woman &amp; it'd be a 1st just as bad as those who voted for Ob https://t.co/sNHv6CydII
RobynTebo_|musicnews_facts|0.0|0.0|1.0|0.0|RT @musicnews_facts: Rihanna wearing a shirt of a picture of herself wearing a Hillary Clinton shirt. She's with HER! #ElectionDay https://
RobynTebo_||0.0|0.0|1.0|0.0|RT @musicnews_facts: Rihanna wearing a shirt of a picture of herself wearing a Hillary Clinton shirt. She's with HER! #ElectionDay https://
ericd111|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
ericd111|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
MitchGhouse|WesVengeance7|0.296|0.0|0.891|0.109|RT @WesVengeance7: The joke is on Hillary if she wins.She'll have to sit at the desk Monica sat under.
LyndaJoHunt|jaynordlinger|0.4291|0.049|0.832|0.119|RT @jaynordlinger: Dear GOP: Of all elections to forfeit. The one when HILLARY CLINTON is the Dem nominee? Are you serious? What the ...?
crustyJaureguii|chasemylovex|0.4404|0.0|0.873|0.127|RT @chasemylovex: Y'all better be throwing away these troll ballots after y'all post these pics for RTs and vote for Hillary.
crmorrone|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
crmorrone|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Goodnightma|Morty_Fied|-0.3382|0.151|0.757|0.092|RT @Morty_Fied: Seizure alert! Sick Hillary doesn't quite have her sea legs as seen here in #Philadelphia. @Cernovich @JackPosobiec https:/
Goodnightma||-0.3382|0.151|0.757|0.092|RT @Morty_Fied: Seizure alert! Sick Hillary doesn't quite have her sea legs as seen here in #Philadelphia. @Cernovich @JackPosobiec https:/
Deep_37_2000|GovMikeHuckabee|0.0|0.0|1.0|0.0|"RT @GovMikeHuckabee: State Dept says it takes 5 yrs to review 31,000 Hillary emails. Let Comey do it!  He can review 650,000 in 1 week!  ht"
YourstrulyBey|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
PrimaveraCraig|FIirtationship|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
PrimaveraCraig|twitter|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
lizabethdevon|KendrialWtf|0.34|0.0|0.893|0.107|"@KendrialWtf she wants hillary to win but she still noticed that people bashed trump for saying ""hell"" in front of children"
_HeartOfaHustla|ClarenceJWhite|0.0|0.069|0.863|0.069|RT @ClarenceJWhite: I feel like Trump &amp; Hillary are two divorced parents fighting over custody of us but we kinda just wanna go live with g
WearKatelyn|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
daddyhaj|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
BriaEWilliams|pettyblackgirI|-0.7269|0.243|0.757|0.0|RT @pettyblackgirI: Hillary is also racist. Hillary is married to a r*pist. Hillary funds genocide &amp; ethnic cleansing. Quit trying to guilt
vic71208|Madonna|0.8877|0.0|0.605|0.395|RT @Madonna: Last night was. Amazing!!! Save this Country please!!  Vote for Hillary Clinton!  Today is the Day!  https://t
vic71208||0.8877|0.0|0.605|0.395|RT @Madonna: Last night was. Amazing!!! Save this Country please!!  Vote for Hillary Clinton!  Today is the Day!  https://t
NessaaRobles|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
NessaaRobles|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
DMashak|ProfessorF|0.8225|0.0|0.703|0.297|"RT @ProfessorF: Wow another example of Hillary's ""superior"" ground game. That's brilliant. Having election officials tell people who to vot"
48Glo|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
ffukesteban|HausOfBitchs|0.6908|0.0|0.808|0.192|RT @HausOfBitchs: If Hillary wins she must make telephone part 2 happen once she has Gaga and Bey on her side. This is the only chance we h
thullcat|giguerja|-0.4215|0.135|0.865|0.0|"RT @giguerja: This worries me. If Rove also comes out as bullish on Hillary, run for the hills. https://t.co/lTy8mrbXX0"
thullcat|twitter|-0.4215|0.135|0.865|0.0|"RT @giguerja: This worries me. If Rove also comes out as bullish on Hillary, run for the hills. https://t.co/lTy8mrbXX0"
LynnMoo36681123|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
LynnMoo36681123|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
PARRIGARA|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
PARRIGARA|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
miamiartblog|instagram|0.0|0.0|1.0|0.0|ONCE AGAIN! HILLARY CLINTON EVERYONE... MIAMI DADE COLLEGE!!! At Miami Dade College! https://t.co/yascaesSle
ColeStuckey1|KellyTkelly6974|0.0|0.0|1.0|0.0|RT @KellyTkelly6974: If Hillary gets elected America is done
ryanduffy_55|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
ryanduffy_55|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
Laurence_Zl|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Laurence_Zl|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
blueebae|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
blueebae|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
ak24474|TeamTrump|0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
ak24474||0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
TRUnderwood7|RealAlexJones|0.836|0.0|0.47|0.53|"RT @RealAlexJones: If @HillaryClinton Wins, Freedom Dies - https://t.co/xX0l6mK2vc  #ElectionNight"
TRUnderwood7|infowars|0.836|0.0|0.47|0.53|"RT @RealAlexJones: If @HillaryClinton Wins, Freedom Dies - https://t.co/xX0l6mK2vc  #ElectionNight"
holmes_hailey00|eeller33|0.5106|0.0|0.879|0.121|RT @eeller33: let's keep this in mind as we go to the polls today:11% of people said they'd trust Hillary in office14% of people believe
Savannahhjoness|Austin_Texas1|0.8294|0.051|0.562|0.387|"RT @Austin_Texas1: If Hillary wins- God is still GodIf Trump wins- God is still GodI may have lost hope in America, but never in God."
nirvanicvibes|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
rachaellippe|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
Boringjaf|Boringjaf|-0.25|0.25|0.75|0.0|@Boringjaf Hillary is actually Trump in disguise.
warrenswords|twitter|0.0|0.0|1.0|0.0|Pup is staying up for election. She's with Hillary. Probably. https://t.co/iQ9n55hiZp
Politolizer|politics|0.0|0.0|1.0|0.0|POLITICO | Even Hillary Clinton 's campaign did the mannequin... https://t.co/f3lml6aQd7 https://t.co/7OEHQB0Cmm
AllyBendecime|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
joymvundura|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
omggbrit|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
omggbrit|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
TWEETY021163|France24_en|0.0|0.0|1.0|0.0|RT @France24_en: #HillaryClinton #USElection2016 Take a look back at Hillary Clinton's biggest headaches during campaign https://t.co/bHGJm
TWEETY021163|t|0.0|0.0|1.0|0.0|RT @France24_en: #HillaryClinton #USElection2016 Take a look back at Hillary Clinton's biggest headaches during campaign https://t.co/bHGJm
maIoufoy|Khanoisseur|0.0772|0.162|0.664|0.174|"RT @Khanoisseur: glorious montage of Trump flipping on every position he's held-Iraq War, Libya, healthcare, amnesty, hillary... https://t."
maIoufoy||0.0772|0.162|0.664|0.174|"RT @Khanoisseur: glorious montage of Trump flipping on every position he's held-Iraq War, Libya, healthcare, amnesty, hillary... https://t."
__BabyKayyy|chasemylovex|-0.3586|0.127|0.873|0.0|"RT @chasemylovex: no, Hillary is not the ""ideal candidate"" but we still gonna vote for her tho... and we'll deal with sis later, ya hear me"
bebebtisam|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
lydialewiis|TeoHalm|0.3182|0.0|0.796|0.204|"RT @TeoHalm: if you're 18, please go and vote hillary."
smilon713|DavidCornDC|0.0|0.0|1.0|0.0|RT @DavidCornDC: Where Hillary Clinton will declare victory or....something else. https://t.co/4b82Lt4UGB
smilon713|twitter|0.0|0.0|1.0|0.0|RT @DavidCornDC: Where Hillary Clinton will declare victory or....something else. https://t.co/4b82Lt4UGB
iceman120|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
liz_houli|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
liz_houli|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
theriseofgomez|agentscullly|-0.2401|0.213|0.633|0.154|RT @agentscullly: I'm not American but honestly scared for u all+the result will have an impact on the whole world so I better wake up to H
Dat_Boi_Bucky|2AFight|0.0|0.0|1.0|0.0|RT @2AFight: Which would you rather see Hillary get?
DRMBYRNES|TheMarkRomano|0.0|0.0|1.0|0.0|RT @TheMarkRomano: Vote Fraud...Votes for Trump switch to Hillary on Pennsylvania voting machines.Source: https://t.co/BE7P6QeKEZ
DRMBYRNES|pittsburgh|0.0|0.0|1.0|0.0|RT @TheMarkRomano: Vote Fraud...Votes for Trump switch to Hillary on Pennsylvania voting machines.Source: https://t.co/BE7P6QeKEZ
momrails|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
thekilljoydani|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
thekilljoydani|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
creminsmom|HillaryIn2016|-0.4003|0.119|0.881|0.0|@HillaryIn2016 If Hillary worked for a bank (any US Company) &amp;  released Confidential Info.... She is fired... Fire Hillary .... Vote Trump!
kentthonlo|wikileaks|-0.3182|0.119|0.881|0.0|RT @wikileaks: New emails reveal Donna Brazille leaked two more debate questions to Hillary Clinton https://t.co/C9flji5x7I More: https:/
kentthonlo|wikileaks|-0.3182|0.119|0.881|0.0|RT @wikileaks: New emails reveal Donna Brazille leaked two more debate questions to Hillary Clinton https://t.co/C9flji5x7I More: https:/
J7Saluki|nypost|-0.3818|0.157|0.843|0.0|RT @nypost: Donald and Hillary weren't the only ones embarrassing themselves this election season https://t.co/LLQTGEgAVV
J7Saluki|twitter|-0.3818|0.157|0.843|0.0|RT @nypost: Donald and Hillary weren't the only ones embarrassing themselves this election season https://t.co/LLQTGEgAVV
RickeyLane14|RickeyLane14|0.0|0.0|1.0|0.0|"RT @RickeyLane14: After a few months of Trump or Hillary in office America gone text Obama and say ""Hey bighead"""
Danielle_eeee|RH1_ERA|0.5994|0.0|0.755|0.245|RT @RH1_ERA: How y'all voting for Bernie and Bernie voting for Hillary.. Lmao
g59riah|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
mikedrion|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
mikedrion|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
AnnaleeGloria|arzE|0.7865|0.0|0.729|0.271|RT @arzE: voting for Hillary doesn't have to be ur longest yeah boy ever. It can be ur shorter yeah boy ever. Just uhh don't waste ur yeah
drewadams_01|Everything_TN|-0.4767|0.193|0.807|0.0|RT @Everything_TN: Fake Hillary fliers found at the Baker Center on UT's campus https://t.co/5PCnsu9398
drewadams_01|twitter|-0.4767|0.193|0.807|0.0|RT @Everything_TN: Fake Hillary fliers found at the Baker Center on UT's campus https://t.co/5PCnsu9398
Rgmedina93|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
Rgmedina93|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
FreeUs551|DrThomasPaul|0.25|0.0|0.92|0.08|RT @DrThomasPaul: #Election2016 is the one where we set our differences aside and do the right thing. #Trump is the last chance for #Americ
jlg718|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: Florida, its Election Day! Polls are open from 7am-7pm. Confirm your polling place now and go vote for Hillary! https:"
HapaGirl2|vnuek|0.2846|0.0|0.918|0.082|"RT @vnuek: In allegory, America as a strong big fish, but if it chooses rotted head (i.e. Hillary) that only means the end - fish rots from"
nathan_mansour|ryanricco813|0.0258|0.0|0.954|0.046|RT @ryanricco813: A vote for Hillary is a vote for Pusha TA vote for Trump is still a vote for Pusha TNo matter what happens Pusha will
wagenfire1|mitchellvii|0.4404|0.0|0.861|0.139|RT @mitchellvii: I'm noticing the exit polls from MSNBC are dramatically better for Hillary than the ones from Fox.
Cxokie|MoniqueAnnalyss|0.6597|0.079|0.683|0.237|RT @MoniqueAnnalyss: I hope Hillary wins and makes a bill that says no person involved in a reality show or business should be allowed to r
mickthehack|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
leighsdavina|twitter|-0.5319|0.267|0.604|0.129|"""I could care less about him or Hillary"" yet they went on a whole ASS rant about Hillary?  https://t.co/4mvIArK5bM"
sciphex|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
sciphex||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
WitnessLaron|NathanZed|0.5267|0.0|0.848|0.152|RT @NathanZed: my 7 year old cousin just now: is Hellen Keller winning me: whatcousin: Hellen Kellerme: Hillary Clinton? cousin: I dont
Snatching_Soles|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
ItsTheVocal|smh|-0.5574|0.167|0.833|0.0|"The @smh live election blog reports one person has died in a shooting near a polling place in Azusa, California https://t.co/JwmLWwog8d"
ItsTheVocal|smh|-0.5574|0.167|0.833|0.0|"The @smh live election blog reports one person has died in a shooting near a polling place in Azusa, California https://t.co/JwmLWwog8d"
gtrburn|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
gtrburn|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
PBurgrealtor|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
PBurgrealtor|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
2figures2|MissLizzyNJ|0.0|0.0|1.0|0.0|"RT @MissLizzyNJ: In light of the recent revelations about #SpiritCooking, Hillary has updated her campaign logo. https://t.co/5xZx2Gafkz"
2figures2|twitter|0.0|0.0|1.0|0.0|"RT @MissLizzyNJ: In light of the recent revelations about #SpiritCooking, Hillary has updated her campaign logo. https://t.co/5xZx2Gafkz"
saveAmerica123|garydurbin2|0.3802|0.0|0.607|0.393|@garydurbin2 Please vote Hillary! https://t.co/7tgyEmAfnb
saveAmerica123|rollingstone|0.3802|0.0|0.607|0.393|@garydurbin2 Please vote Hillary! https://t.co/7tgyEmAfnb
raidersrant|pote_anna|0.4767|0.0|0.763|0.237|@pote_anna @ChandraMJordan @EricTrump show respect to your next president Hillary Clinton
kcsilkey|arzE|0.7865|0.0|0.729|0.271|RT @arzE: voting for Hillary doesn't have to be ur longest yeah boy ever. It can be ur shorter yeah boy ever. Just uhh don't waste ur yeah
jaleel_bee|Beygency|0.6825|0.0|0.797|0.203|"RT @Beygency: It's so true. If she'd voted for Hillary, she would've eaten up the chance to capitalize on white feminism. Snake voted for S"
REB117|realDonaldTrump|0.0258|0.107|0.78|0.112|@realDonaldTrump Hillary telling Bill to make sure the jet has enough gas to go non stop to UAE
Chardnaeee|marwannafuq|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
Chardnaeee|twitter|0.7717|0.0|0.628|0.372|RT @marwannafuq: I hope Hillary Clinton helps black people the way black people are helping her https://t.co/trWnHY7M9J
drunkenpastxls|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
drunkenpastxls|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Ajax2847|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Ajax2847|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
kateloving|HAGOODMANAUTHOR|0.765|0.0|0.763|0.237|RT @HAGOODMANAUTHOR: TRUMP WINS NORTH CAROLINA AND OHIO!!! UH OH... HILLARY BOTS... TRUMPY COMING TO GET YOU!!! #ElectionNight #BernieSande
seanwlknsn|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
LisaPizza9|Politics1516|-0.5754|0.199|0.801|0.0|RT @Politics1516: INSANE! PA Poll Workers Handing Out Instructions How To Vote For Hillary https://t.co/MKsAjewCZ6 https://t.co/60Ei17wrVY
LisaPizza9|newsninja2012|-0.5754|0.199|0.801|0.0|RT @Politics1516: INSANE! PA Poll Workers Handing Out Instructions How To Vote For Hillary https://t.co/MKsAjewCZ6 https://t.co/60Ei17wrVY
bettercallicaro|trumpconcerts|-0.296|0.187|0.696|0.117|RT @trumpconcerts: Bon Jovi. Sounds German. We fought them in wars. Always keep an eye on those people. If Hillary wins we'll all be living
kileyycass|MorrisonKrystan|-0.3182|0.223|0.777|0.0|RT @MorrisonKrystan: Me if Hillary loses the election https://t.co/GUHV8QmZi1
kileyycass|twitter|-0.3182|0.223|0.777|0.0|RT @MorrisonKrystan: Me if Hillary loses the election https://t.co/GUHV8QmZi1
alwaysafriend2|FaithRubPol|-0.5106|0.202|0.798|0.0|RT @FaithRubPol: Hillary: sane person who is socially awkward and imperfect.Trump: madmanBuy a damn history book. Your life could becom
urbangrowthsf|TheMikeLawrence|0.0|0.0|1.0|0.0|RT @TheMikeLawrence: Hillary is going to become the first female president and all she had to do was go up against the human embodiment of
UnicornxGlits|memeprovider|-0.1695|0.196|0.804|0.0|"RT @memeprovider: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
lifeofsab98|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
lifeofsab98|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
BoothRegboo|navyseal6|-0.6808|0.189|0.811|0.0|"RT @navyseal6: You really have to sit back and ask yourself this question, how can anyone vote for Hillary, she lies to you, she lies about"
mmunro91|bononcheeknee|-0.2732|0.141|0.758|0.101|RT @bononcheeknee: For all those saying Hillary will make the world safer: she wants a no-fly zone in Syria and war with nuclear power.
SalouaAmara_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
SalouaAmara_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
MarieHyde|twitter|0.2023|0.124|0.706|0.171|Now let's hope Hillary low information voters don't  believe IT will bring change https://t.co/S9CaPjjzTx
leastimnotu|DVATW|0.5106|0.0|0.87|0.13|RT @DVATW: Bill Clinton tried to cheer up Hillary today by reminding her that Mandela wasn't elected president until after serving 27 yrs i
nicolegerace|JakeRomano3|0.0|0.0|1.0|0.0|RT @JakeRomano3: If you vote Hillary Clinton to be the next president of this country lmk so I can unfollow you
shazuga|WhitestRabbit_|-0.4753|0.208|0.652|0.14|RT @WhitestRabbit_: A vote for Hillary is not actually a vote for Hillary... but for the devil himself.. Vote for Trump to save America!
dhcalalily28|HispanicsTrump|0.6305|0.0|0.803|0.197|RT @HispanicsTrump: Anybody that's still on the fence please think about the future of our country! We can't pass a country ruined by Hilla
pure_jadore|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
pure_jadore|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
TiffinyKC|AFP|0.0|0.0|1.0|0.0|"RT @AFP: A large Hillary for America sign is displayed at the Jacob K. Javits Center in New York, where Clinton's #ElectionNight event is h"
Mfnaughton|Inc|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
Mfnaughton|t|0.3612|0.0|0.872|0.128|RT @Inc: A Nobel Prize-Winning Economist Explains the 1 Thing That Hillary Clinton and Donald Trump Agree On @josephestiglitz https://t.co/
kellybeeeean|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
julieoakman727|K1erry|0.4939|0.0|0.842|0.158|RT @K1erry: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/eKtDR5quR0 via @gatewaypu
julieoakman727|thegatewaypundit|0.4939|0.0|0.842|0.158|RT @K1erry: More Philly Voter Fraud=&gt; Election Workers Hand Out Instructions to Vote Hillary (VIDEO) https://t.co/eKtDR5quR0 via @gatewaypu
quicksi79085962|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
quicksi79085962|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
zayngecko|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Igbtlahey|freckledbutt|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
Igbtlahey|twitter|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
El_Number_Juan1|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
80sRetroPics|nytimes|0.0|0.0|1.0|0.0|#Vintage #Retro #80s How the FBI Reviewed Thousands of Emails in One Week - New York Times https://t.co/cg44qwqLw6
RosieBud521|Scarlett210|-0.6597|0.234|0.766|0.0|RT @Scarlett210: If U can vote 4 #Hillary when you KNOW she's seriously ill maybe U shld forget ur enormous #Obamacare payt &amp; go to the hos
darkblue714|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
UdvTANBgkh9NQth|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
cyrustvdahs|twitter|0.0|0.0|1.0|0.0|Vote Hillary Bitchessssss!!!#ElectionNight https://t.co/2NYEb0dkn0
terriertot|AMTrump4PRES|0.128|0.13|0.722|0.148|RT @AMTrump4PRES: #IAmVotingBecause My dad didn't sacrifice &amp; serve during 2 wars only 2C R great country become part of the #Hillary &amp; #So
PoliticsPeach|missynorris411|0.0|0.117|0.765|0.117|RT @missynorris411: @PoliticsPeach @kurteichenwald @wise_diva Hillary Clinton is a pariah if she loses. How does Obama pardon a foundation?
eye_picard|TarikawiPeace|0.2023|0.108|0.755|0.137|RT @TarikawiPeace: I didn't know Hillary's mother was an orphan abandoned by her parents. What an amazing turn it would be when her daughte
Hundredod_lF|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Hundredod_lF|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
CwbyG2|worldnetdaily|0.0|0.0|1.0|0.0|@worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/RxXiAwbGkW #Texas
CwbyG2|wnd|0.0|0.0|1.0|0.0|@worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/RxXiAwbGkW #Texas
TRUMPNEXTPRES16|nationdivided|-0.7959|0.336|0.664|0.0|RT @nationdivided: Indiana is joining Kentucky saying Hell No to Hillary! Go Trump #MAGA #Election2016 https://t.co/LvElXqBRef
TRUMPNEXTPRES16|twitter|-0.7959|0.336|0.664|0.0|RT @nationdivided: Indiana is joining Kentucky saying Hell No to Hillary! Go Trump #MAGA #Election2016 https://t.co/LvElXqBRef
kat_niicole|RickyRodge|0.0|0.0|1.0|0.0|RT @RickyRodge: Your MCM voted for Hillary 
windshade1|JkgaddisJulie|-0.4184|0.112|0.888|0.0|RT @JkgaddisJulie: RETWEET!! Heard CNN and Fox are colluding and will be calling FL for Hillary prior to all votes being counted. Trying 2
GGNewMusic|GlobalGrind|0.0|0.0|1.0|0.0|RT @GlobalGrind: Let the kids do the talking  #ElectionNight https://t.co/Px9vyA08M7 https://t.co/6jnaYOguj5
GGNewMusic|globalgrind|0.0|0.0|1.0|0.0|RT @GlobalGrind: Let the kids do the talking  #ElectionNight https://t.co/Px9vyA08M7 https://t.co/6jnaYOguj5
TVWithGG|GlobalGrind|0.0|0.0|1.0|0.0|RT @GlobalGrind: Let the kids do the talking  #ElectionNight https://t.co/Px9vyA08M7 https://t.co/6jnaYOguj5
TVWithGG|globalgrind|0.0|0.0|1.0|0.0|RT @GlobalGrind: Let the kids do the talking  #ElectionNight https://t.co/Px9vyA08M7 https://t.co/6jnaYOguj5
LifestyleWithGG|GlobalGrind|0.0|0.0|1.0|0.0|RT @GlobalGrind: Let the kids do the talking  #ElectionNight https://t.co/Px9vyA08M7 https://t.co/6jnaYOguj5
LifestyleWithGG|globalgrind|0.0|0.0|1.0|0.0|RT @GlobalGrind: Let the kids do the talking  #ElectionNight https://t.co/Px9vyA08M7 https://t.co/6jnaYOguj5
57orm|qSTuN|0.7783|0.0|0.469|0.531|@qSTuN do you think hillary is better? lmao
ChaseFischbach|TheOneandOnIyUS|0.7096|0.0|0.753|0.247|RT @TheOneandOnIyUS: The joke is on Hillary if she wins. She'll have to sit at the desk Monica sat under.
crunchrocket|twitter|-0.3182|0.204|0.796|0.0|I just realized Hillary could be part of Ghost Fighter... https://t.co/OsQ9g7gMb0
LemoineDwight|hboulware|0.5719|0.0|0.654|0.346|"@hboulware trump won nom, the saboteurs elected Hillary"
emilee_tolleson|sav_leger|-0.4678|0.179|0.751|0.07|RT @sav_leger: You can't possibly label all Trump supporters racist but get offended when people assume you live off of welfare bc you supp
WyeOtter|ameeritalsham|-0.4215|0.138|0.804|0.058|"RT @ameeritalsham: Hillary Clinton: ""I want the Iranians to know, that if I'm the president, we will attack Iran"" https://t.co/FMb2jIqIRF"
WyeOtter|twitter|-0.4215|0.138|0.804|0.058|"RT @ameeritalsham: Hillary Clinton: ""I want the Iranians to know, that if I'm the president, we will attack Iran"" https://t.co/FMb2jIqIRF"
Juuwah|Ohh_Spazz|-0.8586|0.367|0.568|0.066|"@Ohh_Spazz Hillary is definitely a more qualified political evil but to call her the ""lesser evil"" is kinda meh to me."
EmuCatapults|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
OneLastMyth|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
OneLastMyth|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
MaryElizaMurphy|RihannaReplay|0.5719|0.0|0.519|0.481|RT @RihannaReplay: Hillary won. https://t.co/tuxGpgRlS4
MaryElizaMurphy|twitter|0.5719|0.0|0.519|0.481|RT @RihannaReplay: Hillary won. https://t.co/tuxGpgRlS4
bigbill_ontw|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana 0.6% reporting TRUMP 69.8% | Hillary 26.4%  massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Elect
sambotello2|WeekendSchemers|-0.3818|0.245|0.755|0.0|RT @WeekendSchemers: This is embarrassing. Hillary vs Hillary https://t.co/59K9hRKTe7
sambotello2|twitter|-0.3818|0.245|0.755|0.0|RT @WeekendSchemers: This is embarrassing. Hillary vs Hillary https://t.co/59K9hRKTe7
Aarec_Larsen99|jakegusto|-0.296|0.121|0.879|0.0|"RT @jakegusto: And from that day forth, no child was ever named 'Hillary' or 'Donald' again... #ElectionDay"
changeisneeded_|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
changeisneeded_|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
somekindofdrugg|brendonSkolat|0.0|0.0|1.0|0.0|RT @brendonSkolat: Hillary or Trump could never https://t.co/GMCRutTvNp
somekindofdrugg|twitter|0.0|0.0|1.0|0.0|RT @brendonSkolat: Hillary or Trump could never https://t.co/GMCRutTvNp
CatsandTay|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
CatsandTay|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
Texgalleslie|BocaRatonRC|0.4404|0.0|0.854|0.146|RT @BocaRatonRC: Who better to torch Hillary to a crisp on election eve than firebrand Tomi Lahren? https://t.co/rnfeyqgAOD https://t.co/4Z
Texgalleslie|bizpacreview|0.4404|0.0|0.854|0.146|RT @BocaRatonRC: Who better to torch Hillary to a crisp on election eve than firebrand Tomi Lahren? https://t.co/rnfeyqgAOD https://t.co/4Z
MEdwardsSmart|FoxNews|-0.4767|0.306|0.568|0.127|@FoxNews it's obvious all you morons are for crooked witch hillary. You are no better than CNN
Chimp999|Chimp999|-0.6289|0.228|0.772|0.0|"RT @Chimp999: @cedric_persaud @JamieRJN @WayneDupreeShow SO, YOU AGREER WITH HILLARY THAT ALL AMERICANS ARE STUPID"
angelatherunner|elias_chairez|-0.2348|0.212|0.635|0.153|RT @elias_chairez: People giving Hillary their vote so Trump won't win: https://t.co/0SfLCKj03a
angelatherunner|twitter|-0.2348|0.212|0.635|0.153|RT @elias_chairez: People giving Hillary their vote so Trump won't win: https://t.co/0SfLCKj03a
Lipanantsi|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
bzazzie|TheDonaldNews|-0.68|0.272|0.728|0.0|RT @TheDonaldNews: 62% Of Florida Exit Poll Say Hillary Server Bothered Them Severely! #FoxNews #Hannity #Dobbs https://t.co/LtdbpUP9Qy
bzazzie|twitter|-0.68|0.272|0.728|0.0|RT @TheDonaldNews: 62% Of Florida Exit Poll Say Hillary Server Bothered Them Severely! #FoxNews #Hannity #Dobbs https://t.co/LtdbpUP9Qy
SteadyJalen|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Babylayyyy_|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Wanda11111|JUDAHsCHILDREN|0.7003|0.0|0.746|0.254|"RT @JUDAHsCHILDREN: @mike_58stingray actually true; Hillary wrote her thesis on Marxist Alinsky her mentor&amp; idol, Alinsky dedicated bk Rule"
mommabear405|xebec78|-0.3818|0.157|0.843|0.0|RT @xebec78: Hillary asks for an extension in Durham county NC because she's losing. https://t.co/pAhnyDSXHU
mommabear405|mcclatchydc|-0.3818|0.157|0.843|0.0|RT @xebec78: Hillary asks for an extension in Durham county NC because she's losing. https://t.co/pAhnyDSXHU
zckwilhelm|EmRyannPelt|-0.4767|0.162|0.838|0.0|RT @EmRyannPelt: If you voted for Hillary just because she is a female you're what's wrong with America
StephenBus|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
StephenBus|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
nobscoffeemom|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
nobscoffeemom|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
DanieleDalton|chip_burns|0.5267|0.0|0.825|0.175|@chip_burns @kincannon_show @MagnificentOne_ I used to be. Not so much now. Where is the wisdom in electing Hillary 
MichaelMajor12|kazueger1|0.0|0.0|1.0|0.0|RT @kazueger1: Trey Gowdy Says FBI Investigation Into Hillary Clinton's Emails Isn't Over https://t.co/TUe0i9gZPv
MichaelMajor12|westernjournalism|0.0|0.0|1.0|0.0|RT @kazueger1: Trey Gowdy Says FBI Investigation Into Hillary Clinton's Emails Isn't Over https://t.co/TUe0i9gZPv
dwzd|HillaryClinton|0.0|0.0|1.0|0.0|"RT @HillaryClinton: Ohio, it's Election Day! Polls are open from 6:30am-7:30pm. Confirm your polling place now and go vote for Hillary!  ht"
Farah_Raisi|Palespanish|0.5719|0.0|0.764|0.236|RT @Palespanish: The Middle East if Hillary Clinton wins the election #Election2016 https://t.co/szTeIAKTdF
Farah_Raisi|twitter|0.5719|0.0|0.764|0.236|RT @Palespanish: The Middle East if Hillary Clinton wins the election #Election2016 https://t.co/szTeIAKTdF
The_Uhlexissss|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
KatelynMason11|alexsmith1636|-0.2411|0.109|0.891|0.0|"@alexsmith1636 can you imagine? ""Once again, I am not a fan of Hillary. But once again, I am a democrat.....once again."""
PaulGoodmanCH|Colin_Bloom|0.5719|0.0|0.871|0.129|RT @Colin_Bloom: If #Hillary wins and serves full 4 yrs then there would have been a #Clinton or a #Bush in the West Wing for 36 out of 40
AubreyXOSel|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
AubreyXOSel|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
wolfgang_eric|LeighPatrick|0.0|0.0|1.0|0.0|"RT @LeighPatrick: Given the reports flooding in nationwide, you either vote Hillary or the machine votes Hillary for you. #Corruption #elec"
Sand__Man4|hanstan002|0.0|0.0|1.0|0.0|RT @hanstan002: rt for trumpfav for hillary
AyeeItsBrooke_|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
ForeignnBiii|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ForeignnBiii|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
mms5048|kylegriffin1|0.6369|0.0|0.846|0.154|"RT @kylegriffin1: Clinton camp out w/ new behind-the-scenes vids of HRC, best may be Bill jumping up and down after the 1st debate: https:/"
mms5048||0.6369|0.0|0.846|0.154|"RT @kylegriffin1: Clinton camp out w/ new behind-the-scenes vids of HRC, best may be Bill jumping up and down after the 1st debate: https:/"
isataharmiller|mitchellvii|0.4404|0.0|0.861|0.139|RT @mitchellvii: I'm noticing the exit polls from MSNBC are dramatically better for Hillary than the ones from Fox.
Idntneedtwitta|E_FOST|0.0|0.0|1.0|0.0|RT @E_FOST: Bih Kentucky is 68 Trump 32 Hillary... I don't even need to drive through that state 
ph3ezus|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ph3ezus|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
SicilianGirl208|kincannon_show|0.0|0.0|1.0|0.0|"RT @kincannon_show: Just saw national 2 p.m. exit poll data that's not public. Trump is STOMPING Hillary. Book those tickets to Canada now,"
London_Lady|CleanCutBiz|0.0|0.0|1.0|0.0|RT @CleanCutBiz: Hillary Clinton has a message for  Pantsuit Nation - https://t.co/ssUefVuEFQ #SocialMedia #SocialMarketing https://t.co/Up
London_Lady|mashable|0.0|0.0|1.0|0.0|RT @CleanCutBiz: Hillary Clinton has a message for  Pantsuit Nation - https://t.co/ssUefVuEFQ #SocialMedia #SocialMarketing https://t.co/Up
kttnmutt|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
pmswolfy|AtlTeaPartyLove|0.0|0.0|1.0|0.0|"RT @AtlTeaPartyLove: If your Role Models are Jay Z, Beyonce and GaGa. You voted for Hillary because they told you to. Then, you already los"
wa7csg3|a|0.3612|0.121|0.667|0.212|Optimism From Hillary Clinton and Darkness From Donald Trump at Campaigns End https://t.co/I4Tj9o9Ef8
VictoriaPlowiec|JoeyGraceffaTranslation|0.7964|0.0|0.679|0.321|@JoeyGraceffaTranslation: 57% of Poles believe that Hillary would be a better president than Trump. I love my coun https://t.co/dLa1Iidzor
VictoriaPlowiec|twitter|0.7964|0.0|0.679|0.321|@JoeyGraceffaTranslation: 57% of Poles believe that Hillary would be a better president than Trump. I love my coun https://t.co/dLa1Iidzor
__theRealKarma|twitter|-0.732|0.291|0.709|0.0|Exactly! It's more people to vote for than just Donald or Hillary. People so damn ignorant https://t.co/VMPgwTaYPD
EmilyJauregui96|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
EmilyJauregui96|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
glamourmag|glamour|0.0|0.0|1.0|0.0|WHOA. https://t.co/wFeQ1aDnpr
anne436|mayarajamani|-0.0516|0.113|0.781|0.105|"RT @mayarajamani: Alexandra Imbroscia, 22, is here at Hillary's block party with her mom Nivia Vieva, 62. ""We're here for history,"" Vieva s"
80sRetroPics|usatoday|0.197|0.0|0.887|0.113|#Vintage #Retro #80s Hillary Clinton calls voting for herself a 'most humbling feeling' - USA TODAY https://t.co/9FojUMVVEt
JScruisen|GeorgeHWBush|-0.723|0.302|0.615|0.083|"@GeorgeHWBush It's about the Supreme Court! I didn't like either, but don't want Hillary setting the SC! Very disappointed in the Bush's!"
deeknee_shhaa|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
deeknee_shhaa|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
glazedserenity|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
glazedserenity|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
leezvibes|twitter|0.3612|0.0|0.848|0.152|Us: Hillary you going to do all the stuff you promised us right ?Hillary : https://t.co/AG2E2ZVjue
Diaz__Kevin|ChuBoi|0.5927|0.0|0.778|0.222|RT @ChuBoi: I want to believe it'll be a landslide for Hillary on #electionnight but Brexit makes me think twice lol
CChristophr154|MattMcFarland3|-0.128|0.159|0.701|0.14|@MattMcFarland3 @WFSBnews Likely wait till close to end to know how many dead people to bring in to get Hillary a win.
maxdesl|tluethje|0.4588|0.0|0.84|0.16|"RT @tluethje: Easy vote. I can confidently say Hillary has lead to the deaths of multiple Americans. Trump has a big mouth, but he hasn't k"
elodievogel|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
elodievogel|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
Humanatur3|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Humanatur3|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
dappage5|youtube|-0.6037|0.282|0.718|0.0|DONALD TRUMP'S PRAYER WARRIORS JUST DROPPED A BOMB ON HILLARY CLINTON...... https://t.co/lWgI92Ebp1
VampyDeer948|philsadelphia|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
VampyDeer948|twitter|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
catheriines|freckledbutt|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
catheriines|twitter|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
samavsfan|BarSouthNCelly|0.3612|0.0|0.898|0.102|RT @BarSouthNCelly: Having to vote for Donald Trump or Hillary Clinton is like asking someone to watch Mike Milbury or Pierre McGuire talk
larsencarly|NPR|0.0|0.0|1.0|0.0|RT @NPR: A spokesman for former President George W. Bush confirms to NPR that he and his wife voted for neither Donald Trump nor Hillary Cl
saraemmaanne|ed_hooley|-0.8769|0.404|0.485|0.111|RT @ed_hooley: HILLARY'S VP TIM KAINE REFUSED TO HELP ME. DAUGHTER KILLED BY ILLEGAL IMMIGRANT #ElectionDay #ElectionNight #RAW https://t.
saraemmaanne||-0.8769|0.404|0.485|0.111|RT @ed_hooley: HILLARY'S VP TIM KAINE REFUSED TO HELP ME. DAUGHTER KILLED BY ILLEGAL IMMIGRANT #ElectionDay #ElectionNight #RAW https://t.
joshsmith1805|DavidPlattUKIP|-0.1511|0.067|0.933|0.0|"RT @DavidPlattUKIP: All these polls putting Hillary ahead. The one thing they can't predict is DT's silent vote, the ones that won't admit"
BarrettSammm|PriceParker2|-0.8126|0.346|0.654|0.0|"RT @PriceParker2: If voting for Trump makes you a racist, does voting for Hillary make you a criminal?"
mcchlovin_|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
deannafung|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
deannafung|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
StonedPhillyFan|elctrceye|0.2732|0.129|0.632|0.239|@elctrceye There's going to be a war either way yeah but at least Hillary is competent
MarkBapst1|twitter|0.0|0.0|1.0|0.0|Did they look under Hillary's bed! https://t.co/D4xtC9CR8p
ScholtenJacob|youngdeuey|-0.25|0.25|0.533|0.217|"@youngdeuey @JaydaJolene @2MichaelDunlap3 they're both old, rich and racist. Bad point to rest on for Hillary supporters in my opinion"
Hailey_1190|jamiedupree|0.1779|0.182|0.579|0.24|"@jamiedupree Hillary's supporters have no brain cells, am I right?"
wavvycee|6PAPl|0.4404|0.0|0.879|0.121|RT @6PAPl: if kodak black believes hillary can do a good job with our country then we gotta go vote for hillary https://t.co/RWmwK8wHUR
wavvycee|twitter|0.4404|0.0|0.879|0.121|RT @6PAPl: if kodak black believes hillary can do a good job with our country then we gotta go vote for hillary https://t.co/RWmwK8wHUR
SwiftieMahomie|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
Josheezy_|BarSouthNCelly|0.3612|0.0|0.898|0.102|RT @BarSouthNCelly: Having to vote for Donald Trump or Hillary Clinton is like asking someone to watch Mike Milbury or Pierre McGuire talk
troijohnna|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
troijohnna|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
FirebaughNorman|co_firing_line|0.5267|0.0|0.764|0.236|"OPINION: If Trump Edges Clinton, Will Hillary Go Gracefully? https://t.co/5aH7mgXmEK via @co_firing_line"
FirebaughNorman|conservativefiringline|0.5267|0.0|0.764|0.236|"OPINION: If Trump Edges Clinton, Will Hillary Go Gracefully? https://t.co/5aH7mgXmEK via @co_firing_line"
Blake__Lauren|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Blake__Lauren|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
NimciRdz|imashbuttons|-0.0516|0.134|0.743|0.124|RT @imashbuttons: Why Hillary look like she bout to ask Yugi's grandpa bout some damn cards https://t.co/FZ4H3bLIoK
NimciRdz|twitter|-0.0516|0.134|0.743|0.124|RT @imashbuttons: Why Hillary look like she bout to ask Yugi's grandpa bout some damn cards https://t.co/FZ4H3bLIoK
TheMusicMamaB|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
TheMusicMamaB|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
CarterReed11|awoll2016|0.296|0.0|0.891|0.109|"RT @awoll2016: @AdelleNaz @BreitbartNews Where are Hillary's pop star luciferians singing the National Anthem? Oh yeah, that's right, they"
PearlTommy5|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
PearlTommy5|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
tsmcdonald28|HoltBlack05|-0.4404|0.367|0.633|0.0|RT @HoltBlack05: Hillary Clinton hates puppies
SincerelyQuin_|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
SincerelyQuin_|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Toastiewiththe|TMZ|0.2755|0.0|0.85|0.15|RT @TMZ: Hillary Clinton -- Don't Mess With My Muscle (PHOTO GALLERY) https://t.co/A9vmCznVBk
Toastiewiththe|tmz|0.2755|0.0|0.85|0.15|RT @TMZ: Hillary Clinton -- Don't Mess With My Muscle (PHOTO GALLERY) https://t.co/A9vmCznVBk
boominator|twitter|0.3612|0.173|0.524|0.304|Podesta/Hillary are truly sick individuals supporting Child Trafficking &amp; #SpiritCooking #Occult #ImWithHer https://t.co/O4Wm6Hgi1Y
abiodunsoluade|Nedunaija|0.8126|0.0|0.739|0.261|"RT @Nedunaija: As results start coming in, don't fret if u're for Hillary. The greatest blessing to  Democrats, in my view, is California."
thelifeoftati|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
thelifeoftati|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
favoriterecord||-0.4871|0.193|0.704|0.103|also @ people just voting for trump bc u hate hillary ?????? that's like picking flinging yourself off a cliff on purpose
heatstreet|heatst|0.2023|0.0|0.859|0.141|BUSTED: Top media pundits gave money to Clinton (but there's a catch). https://t.co/onKR1Utvag
FOCVS_Trading|BrockDodd|0.7906|0.0|0.65|0.35|"RT @BrockDodd: Assuming Hillary wins, swinging $XIV is literally free money before market close today."
theyfall4liyah|TheWorldOfFunny|0.0|0.0|1.0|0.0|RT @TheWorldOfFunny: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/rYVq0sC4U5
theyfall4liyah|twitter|0.0|0.0|1.0|0.0|RT @TheWorldOfFunny: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/rYVq0sC4U5
rubyred10123|brandonpearse|-0.1027|0.142|0.735|0.123|RT @brandonpearse: Picking between trump and Hillary is like asking if you wanna be shot or stabbed
rosecal7|lex_looper|0.0|0.0|1.0|0.0|"RT @lex_looper: Hillary stole haiti donations, armed ISIS, covered up child trafficking &amp; she gets the black vote because... Beyonc https:"
howardmclainjr|BlackManTrump|-0.5859|0.183|0.817|0.0|RT @BlackManTrump: Miami4Trump: RT 2ALAW: Voter Fraud In PhiladelphiaPush Button One For HillaryPaid For By The Democratic County.#Elec
LaPecosaAnta|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
LaPecosaAnta|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
gotfamegang|cleanhaylor|0.2118|0.166|0.596|0.238|@cleanhaylor both suck but Hillary is more worth it
BarbaraB777|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
Luxury_etc|teenvogue|0.0|0.0|1.0|0.0|Rihanna Wears a T-Shirt of Herself Wearing a T-Shirt of Hillary Clinton https://t.co/Vlod3PRyyr
twofoneshawty|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
twofoneshawty|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
PureEnergy813|MikePenceVP|-0.7345|0.236|0.764|0.0|RT @MikePenceVP: Hillary's email lies in 45 secondsNo way she should be allowed to serve. Gross &amp; total negligence! #LockHerUp #RT https:
kmfw160|2ALAW|-0.4404|0.231|0.602|0.167|"RT @2ALAW: It's truly a sad day in America when we dismiss all the corruption, voting fraud committed as ""just politics""#Hillary is disqu"
mediohcre|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
mediohcre|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
tanya_vs|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
tanya_vs|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Trump vs Hillary #ElectionDay https://t.co/BRv1x2bYlB
Dezierael|JLaughmiller|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
Dezierael|twitter|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
JoCaseyB|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
ChuckCollier76|kazueger1|0.0|0.0|1.0|0.0|RT @kazueger1: Trey Gowdy Says FBI Investigation Into Hillary Clinton's Emails Isn't Over https://t.co/TUe0i9gZPv
ChuckCollier76|westernjournalism|0.0|0.0|1.0|0.0|RT @kazueger1: Trey Gowdy Says FBI Investigation Into Hillary Clinton's Emails Isn't Over https://t.co/TUe0i9gZPv
Geeeooh15|yvezayntIaurent|-0.5423|0.22|0.78|0.0|"RT @yvezayntIaurent: white person: idk whos worse: hillary or trumplgbtq, women, black people, immigrants, muslims: trump iswhite pers"
cliff_helton24|CloydRivers|0.0|0.0|1.0|0.0|RT @CloydRivers: Im not against a woman bein President. Im just against that woman bein Hillary Clinton. Merica.
sarainestroza8|theScore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
sarainestroza8|thescore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
chloeperkinss|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
audrey_gibbons|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
audrey_gibbons|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
AnnSchm03580293|phil200269|-0.9231|0.489|0.423|0.088|"RT @phil200269: How Is Importing 1Million Syrian Refugee Terrorists and Rapists Going To Help Poverty Stricken Americans, Hillary?#ImVoti"
Alexsmitty_|sassytbh|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
Alexsmitty_|twitter|0.0|0.0|1.0|0.0|RT @sassytbh: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/bqMEchufZd
tritt808|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Babadoosh1|JackPosobiec|0.0|0.0|1.0|0.0|RT @JackPosobiec: Caught! Democrats Campaign for Hillary Inside N Philadelphia Poll https://t.co/FZP07zKb7y
Babadoosh1|periscope|0.0|0.0|1.0|0.0|RT @JackPosobiec: Caught! Democrats Campaign for Hillary Inside N Philadelphia Poll https://t.co/FZP07zKb7y
ThatmustbPharoh|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
ThatmustbPharoh|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
ReidZolinski|TheOneandOnIyUS|0.7096|0.0|0.753|0.247|RT @TheOneandOnIyUS: The joke is on Hillary if she wins. She'll have to sit at the desk Monica sat under.
kyiamonae|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
kyiamonae|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
FreeMilo69|DontTread_2nd|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
FreeMilo69|twitter|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
KareemLumumba|twitter|0.3182|0.0|0.777|0.223|#Trump making sure wifey doesn't vote for #Hillary https://t.co/rU76msyhIc
Kians_Baddie|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
davidprieto08|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
davidprieto08|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
Smedley_Butler|ActualFlatticus|-0.765|0.248|0.752|0.0|RT @ActualFlatticus: Has Hillary Clinton ever said a single word that led you to believe she intends to stop killing people in 7 countries?
Xanthan003|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Xanthan003|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
DebWhit93354460|FoxNews|-0.6449|0.271|0.652|0.077|@FoxNews @HillaryClinton @JakeBGibson She is a criminal! If you want change don't vote Hillary!!!
frazier_ann|kjdrennen|-0.6908|0.322|0.678|0.0|"RT @kjdrennen: .@TheEllenShow whines: @HillaryClinton ""cannot catch a break"" with e-mail scandal https://t.co/EtmQnw681e #TTT16 https://t.c"
frazier_ann|newsbusters|-0.6908|0.322|0.678|0.0|"RT @kjdrennen: .@TheEllenShow whines: @HillaryClinton ""cannot catch a break"" with e-mail scandal https://t.co/EtmQnw681e #TTT16 https://t.c"
GlennManeval|ed_hooley|0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #California #sandiego #OrangeCounty #sacramento #LosAngeles  https://t.
GlennManeval||0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #California #sandiego #OrangeCounty #sacramento #LosAngeles  https://t.
Sparkfoot|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
Sparkfoot|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
jb19tele|rkamienski|0.0|0.0|1.0|0.0|RT @rkamienski: KENTUCKY #exitpollsDonald Trump 66.0%Hillary Clinton 29.8%#ElectionDay
nikemil|kimayad_|0.3612|0.0|0.872|0.128|"RT @kimayad_: Before Hillary Clinton, there was Shirley Chisholm. Thank you for paving the way. #UnboughtAndUnbossed72 #Election2016 http"
HumphryBrokhart|esquire|0.0|0.0|1.0|0.0|Will Ferrell Is Just Your Average Millennial in a New Hillary Clinton Ad - He's with her.  https://t.co/efvfv1i2AO
sophipoo|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
sophipoo|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
Elspeth_Powell|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
Elspeth_Powell|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
bamamom2x|yankeebrit77|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
bamamom2x|twitter|0.0|0.0|1.0|0.0|"RT @yankeebrit77: Why don't these reported ""glitches"" &amp; ""errors"" ever change Hillary votes to Trump? #Rigged #ElectionNight https://t.co/n"
ldrx0|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
ldrx0|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Amyloukingery|FacMagnaAmerica|-0.2023|0.141|0.859|0.0|RT @FacMagnaAmerica: .@JackPosobiec on #Periscope: Hillary Workers Intimidate Voters in Philly https://t.co/MwbHAdq0Zj
Amyloukingery|periscope|-0.2023|0.141|0.859|0.0|RT @FacMagnaAmerica: .@JackPosobiec on #Periscope: Hillary Workers Intimidate Voters in Philly https://t.co/MwbHAdq0Zj
LA_VeryOwn|ItsKrich|-0.7906|0.286|0.714|0.0|RT @ItsKrich: I'm scared of Hillary Clinton because I know exactly what she'll do and I'm scared of Donald Trump because there's no tellin
Wutevuh|TRay1949|0.0|0.0|1.0|0.0|RT @TRay1949: Hillary's Kissin KKK  https://t.co/2RoehKOfht
Wutevuh|twitter|0.0|0.0|1.0|0.0|RT @TRay1949: Hillary's Kissin KKK  https://t.co/2RoehKOfht
JReives04|jozenc|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
JReives04|twitter|0.8625|0.0|0.586|0.414|RT @jozenc: Why Hillary greet all her black friends like she thought they weren't coming to her party? https://t.co/Id0avyHnMZ
__paoeuresti|FIirtationship|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
__paoeuresti|twitter|0.0|0.0|1.0|0.0|RT @FIirtationship: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/LA0LDtKi0P
sardiver3|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
namasteee_|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
hamoudikan|TheSun|0.6204|0.0|0.807|0.193|RT @TheSun: A final poll for the #USElection shows who is most likely to win tonight #USElection https://t.co/6cWAQBvrhi https://t.co/AchWa
hamoudikan|thesun|0.6204|0.0|0.807|0.193|RT @TheSun: A final poll for the #USElection shows who is most likely to win tonight #USElection https://t.co/6cWAQBvrhi https://t.co/AchWa
RushaliSarkar|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
RushaliSarkar|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
twinkIouis|vickto_willy|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
twinkIouis|t|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
cYa_Mahlati|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
cYa_Mahlati|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
HazelOsterhout|PhillyGOP|-0.5859|0.192|0.808|0.0|@PhillyGOP @mshellbeth  Hillary sould be locked uo for commiting fraud thoughout her campaign  #electionday #FoxNews2016  #MAGA #TrashCheats
FenMorgana|gmlively|0.3612|0.0|0.848|0.152|RT @gmlively: I have the Hillary H down pat. These #NastyWomen are ready to #GOTV #ProudToBePA https://t.co/3xvlL7BCQg
FenMorgana|twitter|0.3612|0.0|0.848|0.152|RT @gmlively: I have the Hillary H down pat. These #NastyWomen are ready to #GOTV #ProudToBePA https://t.co/3xvlL7BCQg
tabbyburnsworth|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
F4NZONED|FifaDuaine|0.5719|0.0|0.748|0.252|RT @FifaDuaine: if Hillary wins I'll PayPal everyone $100 that RTs this
JamoneHill|Ma_Ya_Business|-0.5106|0.13|0.87|0.0|RT @Ma_Ya_Business: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY B
hildur789|BreitbartNews|0.4019|0.0|0.597|0.403|RT @BreitbartNews: Special snowflake. https://t.co/k94ncGgmn3
hildur789|breitbart|0.4019|0.0|0.597|0.403|RT @BreitbartNews: Special snowflake. https://t.co/k94ncGgmn3
luispecialone|twitter|-0.2023|0.107|0.893|0.0|There will never be elections in the World as controversial as #Hillary and #Trump   #ElectionNight https://t.co/7OL2bVCLAa
bethvictoire|YUNGMUERTE|0.6369|0.0|0.802|0.198|RT @YUNGMUERTE: I'm gonna try n sleep Hopefully Hillary is president tomorrow morning or maybe someone cooler like snoop dogg and vp is Ma
Sansonel0|musicnews_facts|0.4404|0.0|0.873|0.127|"RT @musicnews_facts: Trump supporters are calling out Hillary Clinton and Lady Gaga for wearing this ""Nazi Hitler"" uniform... When it's Mic"
EricShapiro3|BritsForHill|0.2323|0.101|0.759|0.14|RT @BritsForHill: PLEASE don't assume #Hillary victory is guaranteed...we made that mistake with Brexit. Go out and TAKE IT! #nevertrump
Alyssa_trapani|chanelpuke|-0.1695|0.196|0.804|0.0|"RT @chanelpuke: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
belleponine|taylortetreau|0.5574|0.0|0.816|0.184|RT @taylortetreau: Why is this screenshot from a Hillary campaign video the funniest thing I've ever seen https://t.co/21FbTs3kHb
belleponine|twitter|0.5574|0.0|0.816|0.184|RT @taylortetreau: Why is this screenshot from a Hillary campaign video the funniest thing I've ever seen https://t.co/21FbTs3kHb
capesquad|paul7177|-0.2732|0.231|0.769|0.0|@paul7177 @megynkelly @IngrahamAngle  You're biased according to: https://t.co/q70BVkKich
capesquad|politifact|-0.2732|0.231|0.769|0.0|@paul7177 @megynkelly @IngrahamAngle  You're biased according to: https://t.co/q70BVkKich
cademcfadden|galen_howell|-0.6486|0.515|0.485|0.0|@galen_howell my gun voted for Hillary. :(
nycmidtown|twitter|-0.3875|0.193|0.807|0.0|.#Trump show some respectThe #AmericanFlag is not a hand towel#ElectionNight #ImWithHer #Hillary https://t.co/9wu96oRYK6
slaytina_turner|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
BO3ZBANDENG|twitter|0.6124|0.0|0.688|0.313|Please tell me this is the actual Hillary it would be hilarious https://t.co/gVo8nJfguE
davidgeer11|DrMartyFox|-0.3612|0.189|0.683|0.129|RT @DrMartyFox: #ImVotingBecause We Must Save Babies From #Hillary &amp; #PlannedParenthood Who Will Kill A Baby Minutes Before Birth &amp; S
sweetviolets1|esqonfire|0.357|0.049|0.843|0.108|RT @esqonfire: I wouldn't want failing to vote against Hillary on my conscience &amp; you won't either so GO VOTE TRUMP #MAGA #ElectionDay #Ele
EuanJ_Thomas|Fusion|-0.7351|0.237|0.763|0.0|"RT @Fusion: ""Where are you? Injustice is here.""On the eve of the election, Native Americans fighting for #NoDAPL have a message for Hilla"
ShawtiBroCuz_|youtube|-0.8074|0.422|0.578|0.0|"Tariq Nasheed: Black People Fear Trump's Racism, But Hillary Isn't Different  https://t.co/6ZpGd5XIYq"
tjengland01|MarkDice|-0.4738|0.118|0.882|0.0|RT @MarkDice: Do Hillary voters have to fill out their ballots in blood?  Vote for Trump and let's send that witch into retirement!! #Elect
ManOnTheMoonPGH|bawbbyspears|0.4404|0.0|0.674|0.326|RT @bawbbyspears: Hillary Clinton: *breathes*Trump supporters: https://t.co/UR1h1Gl9DM
ManOnTheMoonPGH|twitter|0.4404|0.0|0.674|0.326|RT @bawbbyspears: Hillary Clinton: *breathes*Trump supporters: https://t.co/UR1h1Gl9DM
cb55uic|shelliecorreia|0.4926|0.0|0.738|0.262|"RT @shelliecorreia: She looks better, and younger, than Hillary! https://t.co/aKPygVOsGL"
cb55uic|twitter|0.4926|0.0|0.738|0.262|"RT @shelliecorreia: She looks better, and younger, than Hillary! https://t.co/aKPygVOsGL"
vylancex|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
vylancex|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
SosaChamberIain|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
Politolizer|politics|0.0|0.0|1.0|0.0|Breitbart | The head of the DNC helped Hillary Clinton... https://t.co/RcyqejvDF4 https://t.co/5ZjJMBEy4H
whyaffiliate|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
Menley897||-0.296|0.215|0.64|0.145|Whether you hate Trump or Hillary@ at least we ALL can agree: https://t.co/h1kBYOb2yW
Menley897|twitter|-0.296|0.215|0.64|0.145|Whether you hate Trump or Hillary@ at least we ALL can agree: https://t.co/h1kBYOb2yW
Itslaurennnnn_|KaneZipperman|-0.6067|0.223|0.722|0.055|"RT @KaneZipperman: we don't care about Trump, we don't care about Hillary, we just want Cory back in the house"
bbrie_|__JonathanJay|-0.6083|0.212|0.698|0.09|RT @__JonathanJay: me: hey how are you doingrandom people: trump is a racist and Hillary is a criminal!!!!!!!!!!!!!!! me: oh ok.
Anon_LosAngeles|FrankLuntz|0.6369|0.0|0.733|0.267|"RT @FrankLuntz: The numbers I'm getting now suggest a nationwide turnout that strongly favors Hillary.And if Hillary does well, so will d"
jayachanel00|jiujiuyulin|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
jayachanel00|twitter|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
_KingYdarb|BasebalIy|0.0|0.0|1.0|0.0|RT @BasebalIy: Hillary bunts
Sck2StOmIck|TrumpTrainNewss|-0.3382|0.123|0.877|0.0|"RT @TrumpTrainNewss: While The Polls are Still Open, FBI Agents Drop the Biggest BOMBSHELL on HILLARY! https://t.co/NTLOjeIUeo https://t.co"
Sck2StOmIck|everynewshere|-0.3382|0.123|0.877|0.0|"RT @TrumpTrainNewss: While The Polls are Still Open, FBI Agents Drop the Biggest BOMBSHELL on HILLARY! https://t.co/NTLOjeIUeo https://t.co"
DmcpartlDavid|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @MaddieAndMichi @enjoynChi @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE
ranpaq|Stonewall_77|0.4847|0.0|0.851|0.149|"RT @Stonewall_77: If This Isn't Torture, What is?THIS is what Hillary Clinton explicitly defended at the third presidential debate."
alyssanbarnette|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
celina_bruner|twitter|0.5719|0.0|0.575|0.425|If they announce Hillary wins https://t.co/9kPFjpjekx
TakeAJillPilll|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
TakeAJillPilll|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
clarisalbr|AprilHayes_|-0.4724|0.139|0.861|0.0|RT @AprilHayes_: Stay in line West Coast!No to Hillary in the Primary! No in the General!#ElectionNight #Election2016 #iVoted #MAGAx3 #Ji
mauxf_|aldairmaruz|0.5719|0.0|0.778|0.222|"RT @aldairmaruz: if Hillary wins, i'll buy everybody who RTs this tacos and horchata."
_brandonsantoyo|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
_brandonsantoyo|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
charprat44|JaredWyand|-0.742|0.285|0.642|0.073|"RT @JaredWyand: Don't be nervous America. We're only facing economic collapse, anarchy, and inevitable civil war if Hillary wins#Election"
BTeboe|INTJutsu|-0.5411|0.143|0.857|0.0|RT @INTJutsu: Hillary destroyed evidence after she received a subpoena to turn over all emails.  She should be in jail for that alone!#Ele
jearuiz|DrMartyFox|-0.3612|0.189|0.683|0.129|RT @DrMartyFox: #ImVotingBecause We Must Save Babies From #Hillary &amp; #PlannedParenthood Who Will Kill A Baby Minutes Before Birth &amp; S
sharlinsky|Liberienne|0.34|0.112|0.68|0.208|RT @Liberienne: Y'all ready for Bill Clinton to be the first lady? Hopefully Hillary cheats on him while in office.
tyramaniece|teenremark|-0.1695|0.196|0.804|0.0|"RT @teenremark: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
diabadassss|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
diabadassss|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
MaggieMay2495|video|0.7701|0.0|0.622|0.378|"Well Said!!! #ElectionFinalThoughts #Election2016  Sean Hannity: If Hillary wins, you own it https://t.co/QHAmNkVA0X"
REALpugner|mtracey|0.4019|0.0|0.906|0.094|"RT @mtracey: Did you know? Lena Dunham is not registered with any party in NY, so therefore could not have voted for Hillary in the NY prim"
graciee_gilbert|Mendevin_|-0.3182|0.315|0.685|0.0|RT @Mendevin_: Hillary Clinton Lost https://t.co/2dVJ5lYQ9g
graciee_gilbert|twitter|-0.3182|0.315|0.685|0.0|RT @Mendevin_: Hillary Clinton Lost https://t.co/2dVJ5lYQ9g
Maxwell_Rei|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Choosing between Trump and Hillary #ElectionDay #myvote2016 https://t.co/JrPa4gKJBj
Maxwell_Rei|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Choosing between Trump and Hillary #ElectionDay #myvote2016 https://t.co/JrPa4gKJBj
ranpogawa|annalevinsonxx|-0.7739|0.226|0.774|0.0|"RT @annalevinsonxx: Im TIRED of this ""crooked Hillary"" rhetoric do u know how many times Donald has broken the law let GO of ur misogynY ht"
boylemansion|aristotiIes|0.0|0.0|1.0|0.0|RT @aristotiIes: election 2016bad end: donald trumpneutral end: jill steingolden end: bernie sanderstrue end: hillary clintonsecret en
sarah_russell00|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
sarah_russell00|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
mattiOgreen|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
mattiOgreen|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
BrodyMorrow20|0997Raaaaquel|0.6239|0.11|0.601|0.29|"RT @0997Raaaaquel: if Hillary wins and makes America shi**y, y'all better not start complaining and crying bc y'all should've voted TRUMP T"
startupjob124|nytimes|0.0|0.0|1.0|0.0|How the FBI Reviewed Thousands of Emails in One Week - New York Times https://t.co/uW0xB7Hts1
guyxxxtrujillo|Michael_4O8|-0.5423|0.226|0.774|0.0|RT @Michael_4O8: fuck Donald trump and Hillary Clinton  ima just move  to Hawaii 
mattfahey_17|NRich_5|0.0258|0.105|0.787|0.109|"RT @NRich_5: If Hillary Clinton takes an early lead tomorrow nobody stress out, its just the Trump supporters haven't got off work yet"
LindaLouJones13|dmon4ever|0.0|0.0|1.0|0.0|RT @dmon4ever:  PODESTA UNCHAINED:#HILLARY?CRONYISM FOREIGN GOVT'Shttps://t.co/7k87SrtzIm#DrainTheSwamp#ElectionDay#myvote2016
toroyyoo|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
toroyyoo|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
J_LadaliaDFI|theScore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
J_LadaliaDFI|thescore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
CharleyAustin|youtube|-0.6037|0.282|0.718|0.0|DONALD TRUMP'S PRAYER WARRIORS JUST DROPPED A BOMB ON HILLARY CLINTON...... https://t.co/POciJlO8XY
sorryimfreddie|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
PoetikPoeta|3_14159265xPi|0.3716|0.0|0.836|0.164|@3_14159265xPi I don't think Hillary is a great candidate either but Trump is a bigot and a half
YouTubeSamLags|fouseyTUBE|0.3036|0.114|0.687|0.199|@fouseyTUBE I'm not surprised that Fousey Tube supporters are voting for Hillary
zoombouse|PixlProphet|-0.7284|0.339|0.661|0.0|RT @PixlProphet: @NC5_JasonLamb @mitchellvii @NC5 So WTF is Hillary even a contender!?
bjonesbrazil|WeNeedTrump|0.0|0.0|1.0|0.0|RT @WeNeedTrump: Twitter wants Donald Trump. 264K retweets for Donald Trump. 35.6K retweets for Hillary Clinton. #MakeAmericaGreatAgain htt
christinaxxxooo|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
LeeMcVeigh|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
mamacato57|NewtTrump|-0.7269|0.316|0.575|0.109|RT @NewtTrump: RETWEET THIS LIKE CRAZY: Hillary's guilty of 70-100 violations of the US Constitution's Emoluments Clause and the media refu
GIANT918|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
GIANT918|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
AgelinaaPaulina|PopCrave|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
AgelinaaPaulina|twitter|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
vliz3|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
vliz3|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
phoenixyvonneee|abbisprong|-0.3182|0.315|0.685|0.0|"RT @abbisprong: ""Hillary Clinton lost"" https://t.co/U95VhqUoDb"
phoenixyvonneee|twitter|-0.3182|0.315|0.685|0.0|"RT @abbisprong: ""Hillary Clinton lost"" https://t.co/U95VhqUoDb"
LenahanChris|weknowwhatsbest|0.5859|0.0|0.847|0.153|"RT @weknowwhatsbest: Should Hillary win, the first item marked on her calendar is to revisit the black community exactly 4 years from now f"
Diamondrosegrfx|surfermom77|0.0|0.0|1.0|0.0|"RT @surfermom77: For 30Yrs. I, Hillary Clinton Have Achieved Every Method of Corruption &amp;Cheated Bernie 2 Be The Democratic Nominee.NOW I'"
politicallyrich|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
politicallyrich|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
SteezyNeesh|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
SteezyNeesh|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ligayarain_|landry_kameron|0.0|0.0|1.0|0.0|RT @landry_kameron: Hillary voters will be in the lead with the polls all morning because republicans have to get off work before they can
Williams_94x|ltsDonaIdTrump_|0.0|0.0|1.0|0.0|RT @ltsDonaIdTrump_: Hillary Clinton's da sells avon
TVnPolitics|freckledbutt|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
TVnPolitics|twitter|-0.2732|0.189|0.699|0.112|RT @freckledbutt: I just got real damn emotional over hillary's suits y'all https://t.co/PTgVxZyTyD
Angiema23Mata|JoeyGraceffa|0.0|0.0|1.0|0.0|@JoeyGraceffa I'm with her HILLARY
racheIschmidt|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
racheIschmidt|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
ambernt19|BigNik|0.7184|0.0|0.682|0.318|RT @BigNik: Hillary Clinton and her crew really did the mannequin challenge this election is such a joke lmfao
startupjob124|usatoday|0.197|0.0|0.861|0.139|Hillary Clinton calls voting for herself a 'most humbling feeling' - USA TODAY https://t.co/lcZvy8G2mU
ohnoitsceleste|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
ohnoitsceleste|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
Damnits_HANNAH|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Damnits_HANNAH|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
fucksolos|melaninrise|0.5719|0.0|0.821|0.179|RT @melaninrise: if Trump  or Hillary  Wins The Election I Am Moving  Out Of The Country  Goodbye America  Hello  U
Kingwoman|BernieSanders|0.4215|0.0|0.865|0.135|RT @BernieSanders: #ImVotingBecause Hillary Clinton will nominate justices who will overturn Citizens United and take back our democracy fr
sheilamterry1|TeamTrump|0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
sheilamterry1||0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
Badgal_stella|RH1_ERA|0.5994|0.0|0.755|0.245|RT @RH1_ERA: How y'all voting for Bernie and Bernie voting for Hillary.. Lmao
movingpart|twitter|-0.6096|0.166|0.834|0.0|it's because they're all catholic so they hate hillary for being pro gay marriage and pro choice that's it literall https://t.co/eKZZqhklCx
courtneyfwagner|twitter|0.0|0.0|1.0|0.0|"Today, I voted for Hillary and then went to a waterfall. #PNW #MadamePresident #ElectionDay https://t.co/PgQlB0IHnC"
popsacuna|CNN|0.0|0.0|1.0|0.0|@CNN @HillaryClinton @realDonaldTrump I will never watch Clinton News Network (cnn) ever again!!! They just as Crooked as Hillary #MAGA
haydalekzandr4L|marimanic216|0.5319|0.0|0.853|0.147|"RT @marimanic216: FOR ANYONE TALKING ABOUT HOW HILLARY DIDN'T SUPPORT THE LGBTQ+: STFU. THAT WAS YEARS AGO. PEOPLE CHANGE, THEIR OPINIONS C"
0DESTOSLEEP|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
0DESTOSLEEP|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
AllenAdkins2|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
tylerbarrett801|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
celina_perez6|iamwill|0.0|0.0|1.0|0.0|RT @iamwill: I voted for Hillary today &amp; I while I was voting I was listening &amp; vibing out to .@AndersonPaak... #votesANDvibes https://t.co
celina_perez6|t|0.0|0.0|1.0|0.0|RT @iamwill: I voted for Hillary today &amp; I while I was voting I was listening &amp; vibing out to .@AndersonPaak... #votesANDvibes https://t.co
mynamehailey|mefeater|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
mynamehailey|twitter|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
la_kil|Ian56789|-0.4767|0.147|0.853|0.0|"RT @Ian56789: NATO is readying 300,000 troops to attack Russia, should Hillary be installed in the White House https://t.co/mfrqJ52xgm"
la_kil|theduran|-0.4767|0.147|0.853|0.0|"RT @Ian56789: NATO is readying 300,000 troops to attack Russia, should Hillary be installed in the White House https://t.co/mfrqJ52xgm"
JoyMulalo|DailyMail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
JoyMulalo|dailymail|0.0|0.0|1.0|0.0|RT @DailyMail: With 1.54% reporting in Kentucky:  Trump 68%  Hillary 28%https://t.co/GMVxvJS7cN #ElectionNight
tsmcdonald28|HoltBlack05|0.0|0.0|1.0|0.0|RT @HoltBlack05: Hillary Clinton wears socks and sandals
DevinVaughAn5|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
DevinVaughAn5|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
Ramsey2222|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Ramsey2222|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
BlakeCole_14|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
BlakeCole_14|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
Truckwreck54|JoeHNewYork|-0.7121|0.248|0.752|0.0|RT @JoeHNewYork: I think #Hillary threw a vase at her pervert husbands head #ElectionNight because he didn't save her a seat to #OrgyIsland
tooshort__|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
aunye__|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
aunye__|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
aIeynamarie|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
aIeynamarie|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
TheMinishKappa|oranvul|0.0|0.0|1.0|0.0|RT @oranvul: Hillary just got my vote https://t.co/btQVZPyR9M
TheMinishKappa|twitter|0.0|0.0|1.0|0.0|RT @oranvul: Hillary just got my vote https://t.co/btQVZPyR9M
RarerThanNiggas|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
RarerThanNiggas|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
CherylLochhead|INTJutsu|-0.5411|0.143|0.857|0.0|RT @INTJutsu: Hillary destroyed evidence after she received a subpoena to turn over all emails.  She should be in jail for that alone!#Ele
_xoae|ComedyWorIdStar|0.0|0.0|1.0|0.0|RT @ComedyWorIdStar: katy Perry dressed as Hillary Clinton. She has zero chill  https://t.co/dDY4yT6qpx
_xoae|twitter|0.0|0.0|1.0|0.0|RT @ComedyWorIdStar: katy Perry dressed as Hillary Clinton. She has zero chill  https://t.co/dDY4yT6qpx
henriqueafm|Goncalo_Hazard|0.0772|0.0|0.794|0.206|RT @Goncalo_Hazard: -Trump e Hillary-Manequim Challenge https://t.co/I22YjpwLLd
henriqueafm|twitter|0.0772|0.0|0.794|0.206|RT @Goncalo_Hazard: -Trump e Hillary-Manequim Challenge https://t.co/I22YjpwLLd
LeeBrocklebank|Bosox3|0.0516|0.138|0.714|0.148|RT @Bosox3: Hillary supporters are blind to the facts that she isn't the right choice #ElectionNight
TyWavy_|6PAPl|0.4404|0.0|0.879|0.121|RT @6PAPl: if kodak black believes hillary can do a good job with our country then we gotta go vote for hillary https://t.co/RWmwK8wHUR
TyWavy_|twitter|0.4404|0.0|0.879|0.121|RT @6PAPl: if kodak black believes hillary can do a good job with our country then we gotta go vote for hillary https://t.co/RWmwK8wHUR
AmericanPat1981|larryelder|0.5859|0.0|0.826|0.174|"@larryelder Trump essentially ran against GOP, Pres Clinton, Pres Obama, Hillary, and media-most qualified candidate ever-should win by 30"
remzelk1|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @ScottBaio @saskamare @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE NEW P
JEL317|bmangh|-0.1531|0.078|0.922|0.0|RT @bmangh: Pregnant woman votes for Hillary Clinton while in labour after stopping at polls en route to hospital https://t.co/Q47PkbqN0j @
JEL317|telegraph|-0.1531|0.078|0.922|0.0|RT @bmangh: Pregnant woman votes for Hillary Clinton while in labour after stopping at polls en route to hospital https://t.co/Q47PkbqN0j @
safahthesafari|Brown_Saraah|0.0|0.0|1.0|0.0|"RT @Brown_Saraah: People saying Hillary is corrupt don't realize that literally ANYWHERE there's lots of money and/or politics involved, th"
ImAlwaysCoolest|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
Your__Highness_|Lexual__|0.3182|0.0|0.905|0.095|RT @Lexual__: Another comment: all the things y'all mentioned Hillary doing I'm sure Trump would have done if he had a career in politics.
JoshCohenRadio|twitter|0.0|0.0|1.0|0.0|Donald Trump and Hillary Clinton will watch the election results tonight from buildings exactly 450 feet apart. Awk https://t.co/56JcLt2tUT
onlystacee|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
onlystacee|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
HomelessQuatchi|TMZ|0.2755|0.0|0.85|0.15|RT @TMZ: Hillary Clinton -- Don't Mess With My Muscle (PHOTO GALLERY) https://t.co/A9vmCznVBk
HomelessQuatchi|tmz|0.2755|0.0|0.85|0.15|RT @TMZ: Hillary Clinton -- Don't Mess With My Muscle (PHOTO GALLERY) https://t.co/A9vmCznVBk
sirenish_19|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
RoseMaryTBA|GovMikeHuckabee|0.0|0.0|1.0|0.0|"RT @GovMikeHuckabee: State Dept says it takes 5 yrs to review 31,000 Hillary emails. Let Comey do it!  He can review 650,000 in 1 week!  ht"
SiCarswell|irishtimes|0.0|0.0|1.0|0.0|Polls closing in GOP-leaning Georgia &amp; Democratic-leaning Virginia shortly: here's feature I did on Georgia:https://t.co/m5425cODhU
shyanne2017_|Parkerdyro_|0.3612|0.0|0.872|0.128|"RT @Parkerdyro_: Voting for Hillary because she is a woman is like considering marching band a sport because they're a ""team"""
lnick2934|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
lnick2934|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
nadjlaa6731|ParksAndRecPics|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
nadjlaa6731|twitter|0.0|0.0|1.0|0.0|RT @ParksAndRecPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/1kSRUaxGAw
Garrett_Downs_|TheWizKhalifa|-0.9022|0.41|0.59|0.0|RT @TheWizKhalifa: People hate Trump because the media made them hate Trump.People hate Hillary because they are paying attention.#Elec
HapaGirl2|RealAlexJones|0.836|0.0|0.47|0.53|"RT @RealAlexJones: If @HillaryClinton Wins, Freedom Dies - https://t.co/xX0l6mK2vc  #ElectionNight"
HapaGirl2|infowars|0.836|0.0|0.47|0.53|"RT @RealAlexJones: If @HillaryClinton Wins, Freedom Dies - https://t.co/xX0l6mK2vc  #ElectionNight"
mintedpotters|polaroidbones|-0.607|0.184|0.816|0.0|RT @polaroidbones: DONT SPLIT THE DEMOCRATIC VOTE TOMORROW CAUSE YOU DONT WANNA BE STUCK HILLARY OR TRUMP! ITS ONLY GONNA LEAVE US WITH TRU
chandlershelzi|JimBurnell|0.5754|0.0|0.747|0.253|RT @JimBurnell: @realDonaldTrump YES BY ELECTING HILLARY CLINTON! And then I unfollow you.
xpload32004|DRUDGE_REPORT|0.3182|0.0|0.827|0.173|RT @DRUDGE_REPORT: Madonna breaks promise to give oral to Hillary voters... https://t.co/obsQ3RlTFO
xpload32004|nydailynews|0.3182|0.0|0.827|0.173|RT @DRUDGE_REPORT: Madonna breaks promise to give oral to Hillary voters... https://t.co/obsQ3RlTFO
buttonlol|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
IMASOONERFAN1|BeladonnaRogers|-0.4019|0.124|0.876|0.0|"RT @BeladonnaRogers: Sen. Tim Kaine, your basic pipsqueak, boycotted PM Netanyahu's address to Congress on #IranDeal. Now he's running with"
deIuxecoldwater|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
Activeviii|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
SGRobinson97|Things4Guys|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
SGRobinson97|twitter|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
DonnaMacfarlane|doublexmag|0.2263|0.121|0.701|0.178|Forget this Hillary is unlikable stuff. Hillary is downright inspiring. https://t.co/M78kmRLSsh via @doublexmag
DonnaMacfarlane|slate|0.2263|0.121|0.701|0.178|Forget this Hillary is unlikable stuff. Hillary is downright inspiring. https://t.co/M78kmRLSsh via @doublexmag
easton_verkamp|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
Kschnappx0|rxphillip|0.5719|0.0|0.829|0.171|RT @rxphillip: If Hillary Clinton wins does that Make Bill Clinton the First Lady or the first nigga or
MaryThrelkeld4|fmlannalisa|0.0516|0.214|0.556|0.23|@fmlannalisa we ask Hillary supporters the same Damn thing.
EmilyCrosley12|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Udyx_|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
AngelaSelina08|CloydRivers|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
AngelaSelina08|amp|0.0|0.0|1.0|0.0|"RT @CloydRivers: To everyone who wants to vote for Hillary just to keep Trump from becomin' President, watch this...https://t.co/TuUpD7Qgcg"
toiletwhore666|gayprincesss|0.8784|0.0|0.674|0.326|RT @gayprincesss: Now is not the time to joke about trump winning. Get up and go vote for Hillary we really cant have a racist prick in off
BelindaSpeight2|Americooligan|0.0|0.0|1.0|0.0|"RT @Americooligan: Trump up 70.5% to Hillary's 25.8% in Indiana. 35,646 votes to 13,049 (1% reporting). #ElectionNight"
Mannix1925|nationdivided|-0.7959|0.336|0.664|0.0|RT @nationdivided: Indiana is joining Kentucky saying Hell No to Hillary! Go Trump #MAGA #Election2016 https://t.co/LvElXqBRef
Mannix1925|twitter|-0.7959|0.336|0.664|0.0|RT @nationdivided: Indiana is joining Kentucky saying Hell No to Hillary! Go Trump #MAGA #Election2016 https://t.co/LvElXqBRef
iamTidus_|WesVengeance7|0.296|0.0|0.891|0.109|RT @WesVengeance7: The joke is on Hillary if she wins.She'll have to sit at the desk Monica sat under.
HaruspexOfHell|Ultraviolet1197|0.0018|0.118|0.763|0.119|"@Ultraviolet1197 Lol, the whole thing is fucking ridiculous and half of these people are voting for Hillary without doing research."
DemBums4Ever|Variety|0.0|0.0|1.0|0.0|RT @Variety: George W. Bush didn't vote for Donald Trump or Hillary Clinton for president https://t.co/JaXKzBWOTY https://t.co/CspXjAF5AS
DemBums4Ever|variety|0.0|0.0|1.0|0.0|RT @Variety: George W. Bush didn't vote for Donald Trump or Hillary Clinton for president https://t.co/JaXKzBWOTY https://t.co/CspXjAF5AS
annaloulively|unsmokabIe|-0.5423|0.22|0.78|0.0|"RT @unsmokabIe: white person: idk whos worse: hillary or trumplgbtq, women, black people, immigrants, muslims: trump iswhite person: i"
LoveeeDommm|Kate_da_Bonbon|-0.2382|0.14|0.86|0.0|RT @Kate_da_Bonbon: They both suck but I'd rather have Hillary as president #ElectionNight
mochabearflex|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
mochabearflex|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
dtotheina|TAXSTONE|0.743|0.0|0.704|0.296|RT @TAXSTONE: I feel like Hillary might win then pull off the mask and still be Donald Trump
prettyakasian|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
prettyakasian|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
adamj_film|TragicAllyHere|0.0|0.0|1.0|0.0|"RT @TragicAllyHere: My 6 yr old: ""They asked at school if I wanted Donald Trump or Hillary Clinton but *tearing up* I don't know, I just wa"
Mountainaires|MeetingEjovwo|0.1655|0.0|0.916|0.084|"@MeetingEjovwo Puerto Ricans, Venezuelans, Colombians, Mexicans in FL for Hillary. Cubans always supported the GOP, but younger Cubans, less"
nancyl367|___RaelynnD___|0.7925|0.0|0.707|0.293|RT @___RaelynnD___: @JuliaSokolowski I am a PROUD transfemale for Trump. Hillary is NOT a friend to #LGBT.She uses groups and causes until
SantyCanolopez|PoeticsNormani|0.7717|0.0|0.309|0.691|RT @PoeticsNormani: Hillary better win
nativeoldcrow|AssangeFreedom|0.2481|0.092|0.761|0.146|RT @AssangeFreedom: @Wikileaks docs proved #Hillary seriously endangered  American security with her private email server! #ImVotingBecause
MazvitaJames|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
MazvitaJames|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
isabelrichardss|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
vipertoxin|youtube|-0.5574|0.286|0.714|0.0|&gt;&gt; Hillary Clinton: Im adamantly against illegal immigrants. - YouTube https://t.co/lCbY2BClf0
Cici0804|RealDonalDrumpf|0.8398|0.0|0.53|0.47|@RealDonalDrumpf @votermolly Wow! A WWII veteran. Congratulations for voting for Hillary Clinton.
GaboooTM|BuzzFeedLGBT|0.4019|0.0|0.828|0.172|RT @BuzzFeedLGBT: People Are Wearing Pantsuits Today To Show Their Support For Clintonhttps://t.co/RjNfsJHwqc https://t.co/oQ0Uc4nBvM
GaboooTM|twitter|0.4019|0.0|0.828|0.172|RT @BuzzFeedLGBT: People Are Wearing Pantsuits Today To Show Their Support For Clintonhttps://t.co/RjNfsJHwqc https://t.co/oQ0Uc4nBvM
glendabelle_11|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
GalInTheGreyHat|KristinHarris|0.7463|0.0|0.71|0.29|RT @KristinHarris: Hillary Clinton left this note in the Pantsuit Nation FB group and now I'll truly never stop crying   https://t.co/bP
GalInTheGreyHat|t|0.7463|0.0|0.71|0.29|RT @KristinHarris: Hillary Clinton left this note in the Pantsuit Nation FB group and now I'll truly never stop crying   https://t.co/bP
croskopi|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
croskopi|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
zachkrzeminski1|lindsaylohan|0.0|0.0|1.0|0.0|RT @lindsaylohan: Heart for Hillary or retweet for Trump!
Dakota_Hays34|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
Purpxpink|bigshitxtalker|0.0|0.0|1.0|0.0|RT @bigshitxtalker: Polls close at 7 pm. Hurry up and get in line and vote for Hillary. https://t.co/rBZu2LjQlJ
Purpxpink|twitter|0.0|0.0|1.0|0.0|RT @bigshitxtalker: Polls close at 7 pm. Hurry up and get in line and vote for Hillary. https://t.co/rBZu2LjQlJ
siaayrom|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
t_spoil|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
t_spoil|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
kingjames104|Stonewall_77|0.4847|0.0|0.851|0.149|"RT @Stonewall_77: If This Isn't Torture, What is?THIS is what Hillary Clinton explicitly defended at the third presidential debate."
chrispkeating|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
chrispkeating|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
miniautomatiste|davidsocomedy's|0.296|0.0|0.891|0.109|Catching up on @davidsocomedy's vids So I can think about something other than Trump or Hillary. It's helping immen https://t.co/t6mtoOwCwu
miniautomatiste|twitter|0.296|0.0|0.891|0.109|Catching up on @davidsocomedy's vids So I can think about something other than Trump or Hillary. It's helping immen https://t.co/t6mtoOwCwu
florbaldassini|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
Shelby_Ryan2125|brittanymacik|0.7506|0.0|0.652|0.348|RT @brittanymacik: All in favor of Texas seceding from the US if Hillary wins
CarverCallie|tedperl|-0.69|0.216|0.784|0.0|@tedperl @DonaldJTrumpJr Nothing works in Haiti when you have #CrookedHillary running it. Look into https://t.co/7Uwqx69GaL Hillary is evil!
CarverCallie|beforeitsnews|-0.69|0.216|0.784|0.0|@tedperl @DonaldJTrumpJr Nothing works in Haiti when you have #CrookedHillary running it. Look into https://t.co/7Uwqx69GaL Hillary is evil!
sonjamart48|Koxinga8|0.7667|0.0|0.662|0.338|RT @Koxinga8: HAPPY ELECTION DAY! FBI Agents Just Surprised Comey With New Hillary Crimes https://t.co/Eafa46JVnq
sonjamart48|angrypatriotmovement|0.7667|0.0|0.662|0.338|RT @Koxinga8: HAPPY ELECTION DAY! FBI Agents Just Surprised Comey With New Hillary Crimes https://t.co/Eafa46JVnq
annhcallaway|HillaryClinton|0.0|0.0|1.0|0.0|@HillaryClinton A Song for you https://t.co/1KW1QsyRiI
annhcallaway|soundcloud|0.0|0.0|1.0|0.0|@HillaryClinton A Song for you https://t.co/1KW1QsyRiI
HolyMindfreak|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
harrysfruitpack|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
American4DJT|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
StephGrobler1|FrankLuntz|-0.6705|0.341|0.537|0.122|@FrankLuntz If you like a corrupt lying sack of shit as #POTUS go for hillary
livfrosty|lilyachty|0.0|0.0|1.0|0.0|RT @lilyachty: Hillary! https://t.co/VZMLR24Y3Y
livfrosty|twitter|0.0|0.0|1.0|0.0|RT @lilyachty: Hillary! https://t.co/VZMLR24Y3Y
mary_mccartney|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
mary_mccartney|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
louiselloyd3|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana 0.6% reporting TRUMP 69.8% | Hillary 26.4%  massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Elect
VoteTrumpPence7|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
OGYoungPrincess|iamdiddy|0.0|0.0|1.0|0.0|hey i voted (for hillary) can i have $500? @iamdiddy
cpalmero27|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
BNB52|shoutout_TAG|0.25|0.0|0.917|0.083|RT @shoutout_TAG: If you live in Florida Ohio Michigan or Pennsylvania you have a chance still to keep Hillary and the establishment out of
partyrt2010|BreitbartNews|0.0|0.0|1.0|0.0|RT @BreitbartNews: Birds of a feather. https://t.co/UdePaJZYyY
partyrt2010|breitbart|0.0|0.0|1.0|0.0|RT @BreitbartNews: Birds of a feather. https://t.co/UdePaJZYyY
The_Uhlexissss|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
kleeoosullivan|1942bs|-0.8304|0.277|0.688|0.034|"RT @1942bs: Black ppl are getting shamed no matter what we choose to do with our vote. We cant win by not voting, voting for Hillary/Trump,"
rns_lake2|Iightmeup|0.0|0.0|1.0|0.0|RT @Iightmeup: Just another reason to vote for Hillary  #ImWithHer https://t.co/djoAYLUs8w
rns_lake2|twitter|0.0|0.0|1.0|0.0|RT @Iightmeup: Just another reason to vote for Hillary  #ImWithHer https://t.co/djoAYLUs8w
Wolffox6|agreatercountry|-0.2481|0.135|0.767|0.099|"RT @agreatercountry: Lying MSM, for the last month is telling us the Latino support was surging for Hillary. CNN Poll shows NOT TRUE!http"
Robbull951|_Makada_|0.8916|0.0|0.608|0.392|"RT @_Makada_: Trump in Manchester, NH: ""Hillary's only allegiance is to herself, her donors, and her special interests! My only special int"
justcallmeKy|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
justcallmeKy|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
pjbowles|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @YoungDems4Trump @enjoynChi @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE
crappers51|CNN|-0.4215|0.135|0.865|0.0|@CNN O I REALLY FEEL FOR HILLARY LETS NOT TALK ABOUT ALL THE LAWS SHE BROKE LETS NOT TALK ABOUT TTTHHHAAAT
jtoufas|BobMacAZ|-0.6908|0.239|0.761|0.0|"RT @BobMacAZ: BREAKING: Hours Before Polls Close, Rape Allegation Sends Hillary Into Tailspin https://t.co/sU3y6q2Bu7 via @USADailyInfo"
jtoufas|dailyinfo|-0.6908|0.239|0.761|0.0|"RT @BobMacAZ: BREAKING: Hours Before Polls Close, Rape Allegation Sends Hillary Into Tailspin https://t.co/sU3y6q2Bu7 via @USADailyInfo"
ranvir01|FrankLuntz|0.6369|0.0|0.733|0.267|"RT @FrankLuntz: The numbers I'm getting now suggest a nationwide turnout that strongly favors Hillary.And if Hillary does well, so will d"
normansreed|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
normansreed|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
rsanterre44|Cory_1077|-0.8159|0.453|0.547|0.0|RT @Cory_1077: #HILLARY WILL BANKRUPT GUN MAKERS BY EXECUTIVE ORDERhttps://t.co/YXWmAZJxND https://t.co/TSLRnmDEMx
rsanterre44|twitter|-0.8159|0.453|0.547|0.0|RT @Cory_1077: #HILLARY WILL BANKRUPT GUN MAKERS BY EXECUTIVE ORDERhttps://t.co/YXWmAZJxND https://t.co/TSLRnmDEMx
trumpquility1|mitchellvii|0.4404|0.0|0.861|0.139|RT @mitchellvii: I'm noticing the exit polls from MSNBC are dramatically better for Hillary than the ones from Fox.
BriannaLeJeunee|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
BriannaLeJeunee|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
dougsmith1946|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
lastname_jeter|JLaughmiller|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
lastname_jeter|twitter|0.4939|0.0|0.714|0.286|RT @JLaughmiller: Hillary vs. Hillary. Pretty eye opening:) https://t.co/7uGMyjsR7j
karenbr01503349|umpire43|0.4019|0.0|0.891|0.109|RT @umpire43: My old Boss Reuters had a poll showing Hillary support nosedived to 36% in last 4 days.They took the poll down a few minutes
L7Feldare|Tehxture|0.0|0.0|1.0|0.0|RT @Tehxture: THESE FUCKING IDIOTS REALIZE TRUMP AND HILLARY ARENT THE ONLY ONES ON THE BALLOT???????????????????
southpaw816|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
LyellBan|BlissTabitha|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
LyellBan|weaselzippers|0.0|0.0|1.0|0.0|RT @BlissTabitha: Freddie Gray Prosecutor Marilyn Mosby Breaks Law By Taking Photo While Voting For Hillary https://t.co/8UcX6CEWcr
TylerC133|OnlineMagazin|-0.5267|0.207|0.714|0.079|RT @OnlineMagazin:  That made my day. Crooked Hillary supporter went into the trap when he wanted to steal the #DonaldTrump shield. ht
CoconutGucci2|porn_horse|-0.7656|0.292|0.708|0.0|RT @porn_horse: Hillary campaigner employed FORBIDDEN MAGIC to do a kickflip in heels. No one is talking about this!!!https://t.co/GD9L0u
CoconutGucci2|t|-0.7656|0.292|0.708|0.0|RT @porn_horse: Hillary campaigner employed FORBIDDEN MAGIC to do a kickflip in heels. No one is talking about this!!!https://t.co/GD9L0u
marcylauren|pablorodas|0.8436|0.0|0.702|0.298|RT @pablorodas: Hillary winning in 7 key states followed by Slate tracker! Great! #tcot #PJNET #GOP #2A #ccot #teaparty #tlot #MAGA #Trump2
_mLr|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
_mLr|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
citzncinematrix|FemMajority|0.0|0.0|1.0|0.0|"RT @FemMajority: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https"
sakurafishguy|twitter|-0.5232|0.214|0.704|0.082|"So the ""hes not winning""  confidence is already out the Hillary supporter window.  Now hes not gonna last his first https://t.co/rRoSj8vTsv"
factanonverba7|marklevinshow|-0.4588|0.333|0.667|0.0|RT @marklevinshow: Disgraced Comey and Lynch https://t.co/dsl7nNuguV
factanonverba7|nationalreview|-0.4588|0.333|0.667|0.0|RT @marklevinshow: Disgraced Comey and Lynch https://t.co/dsl7nNuguV
adelaide_hall3|atensnut|-0.6808|0.167|0.833|0.0|"RT @atensnut: I was 35 years old when Bill Clinton, Ark. Attorney General raped me and Hillary tried to silence me.  I am now 73....it neve"
envydatropic|Treestand_tweet|0.3802|0.0|0.885|0.115|RT @Treestand_tweet: Dude they are still running Hillary commercials give it a break please. I get she didn't use the P word got it!
_whatshername|Jezebel|-0.7269|0.319|0.681|0.0|"RT @Jezebel: All the sad, woke men forced to vote for Hillary Clinton https://t.co/X22INC8Dqa https://t.co/LXAvCNzHX0"
_whatshername|theslot|-0.7269|0.319|0.681|0.0|"RT @Jezebel: All the sad, woke men forced to vote for Hillary Clinton https://t.co/X22INC8Dqa https://t.co/LXAvCNzHX0"
lIbby_annn|UdnSpeak4me|0.0|0.0|1.0|0.0|RT @UdnSpeak4me: Womens rights activists reunite 40 years later to campaign for Hillary Clinton https://t.co/SKC2FlRgp9
lIbby_annn|medium|0.0|0.0|1.0|0.0|RT @UdnSpeak4me: Womens rights activists reunite 40 years later to campaign for Hillary Clinton https://t.co/SKC2FlRgp9
DaddySizzler|jaureologist|-0.0516|0.207|0.591|0.202|RT @jaureologist: I DON'T CARE HOW MUCH Y'ALL HATE BOTH CANDIDATES YOU WILL VOTE FOR HILLARY WHETHER YOU LIKE IT OR NOT I REFUSE TO LET TRU
hanna_felton|twitter|0.0|0.0|1.0|0.0|Go Hillary !! https://t.co/8pFk3ZyaCg
DemiWoehl|talynnsmithh|0.5773|0.0|0.855|0.145|"RT @talynnsmithh: for all u Hillary fans that believe 36 week abortion isn't murder- this is my brother, born @ 28 weeks &amp; i couldn't imagi"
FredSmerlas|worldnetdaily|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
FredSmerlas|wnd|0.0|0.0|1.0|0.0|RT @worldnetdaily: BALLOTS SWITCH TO HILLARY BEFORE VOTERS' EYESObama sends out DOJ monitors to 28 states https://t.co/6RIvNZcoZ2 https:/
SculptNewYork|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
SculptNewYork|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
DerekMiller19|OhioStateDaily|0.0|0.0|1.0|0.0|RT @OhioStateDaily: Donald Trump Hillary Clinton Urban Meyer Urban Meyer 4 President #Election2016 #MyVote2016 https://t.co/r0V2bI7
DerekMiller19|t|0.0|0.0|1.0|0.0|RT @OhioStateDaily: Donald Trump Hillary Clinton Urban Meyer Urban Meyer 4 President #Election2016 #MyVote2016 https://t.co/r0V2bI7
j_queenx|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
j_queenx|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
releeusa|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
teresarc17|mitchellvii|-0.3182|0.206|0.653|0.141|"RT @mitchellvii: If true, this is brutal for Hillary.  She won't match Obama's numbers. https://t.co/z0o069Bv1p"
teresarc17|twitter|-0.3182|0.206|0.653|0.141|"RT @mitchellvii: If true, this is brutal for Hillary.  She won't match Obama's numbers. https://t.co/z0o069Bv1p"
aries1895|GIRLHEFUNNY|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
aries1895|twitter|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
lildg54|BerniedOut|0.5255|0.0|0.834|0.166|"RT @BerniedOut: In Chicago, I had friends waiting last night to vote for 3 hours and moreand we're completely Hillary!"
Just_a_Fiasco|GIRLHEFUNNY|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
Just_a_Fiasco|twitter|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
NOTKASSIE96|RihannaReplay|0.5719|0.0|0.519|0.481|RT @RihannaReplay: Hillary won. https://t.co/tuxGpgRlS4
NOTKASSIE96|twitter|0.5719|0.0|0.519|0.481|RT @RihannaReplay: Hillary won. https://t.co/tuxGpgRlS4
KalaBabu08|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
wldioverbitches|AqueleBlack|0.0|0.0|1.0|0.0|RT @AqueleBlack: Entre o Trump e a Hillary... prefiro o Kanye West...
emilycwalker7|blvckpapii|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
emilycwalker7|twitter|0.0|0.0|1.0|0.0|RT @blvckpapii: Trump vs Hillary at election today  https://t.co/mO8byI0rK1
iammsaraaa|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
iammsaraaa|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
fergesor|StatesPoll|0.0|0.0|1.0|0.0|RT @StatesPoll: Indiana 0.6% reporting TRUMP 69.8% | Hillary 26.4%  massive #TRUMPocrats#TrumpTrain #Maga #VoteTrump #election2016 #Elect
mma_jc|GIRLHEFUNNY|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
mma_jc|twitter|0.5859|0.0|0.703|0.297|RT @GIRLHEFUNNY: If Donald trump or Hillary Clinton win  https://t.co/HxwsonLkP1
TrumpDyke|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
Americans4Gary|Jason4Liberty|0.0|0.0|1.0|0.0|RT @Jason4Liberty: Who are you voting for this #ElectionDay? #NOV8 #Hillary #Trump #GaryJohnson #JillStein #LiveFree #MAGA #ImWithHer #P2 #
lynn5813|OnlineMagazin|-0.5267|0.207|0.714|0.079|RT @OnlineMagazin:  That made my day. Crooked Hillary supporter went into the trap when he wanted to steal the #DonaldTrump shield. ht
rxna21|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
Brookieee1221|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
_mllelbl|AnBressBBC|0.5719|0.067|0.737|0.196|"RT @AnBressBBC: I'm about to walk from the Trump Tower to Hillary's party. Will post about people, supporters or protesters I meet on my wa"
RockyBrown11|hitgirl2now|0.2732|0.0|0.9|0.1|"RT @hitgirl2now: Although Hillary is doing well with white, college educated women, this one voted 4 Trump.  I actually read the Wikileaks"
FatJesusMERZ|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
bradleykarnes|explicitriddle|0.49|0.0|0.757|0.243|@explicitriddle @_PENGUlN don't get me wrong. I know Hillary is gonna win but I don't know why
RobotBrush|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
RobotBrush|thehill|0.0|0.0|1.0|0.0|RT @thehill: Spokesman: George W. Bush did not vote for Clinton https://t.co/AMuzb6nyiM https://t.co/WcqFBXo1YK
Donovanfrom900|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
mlynne3|ed_hooley|0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #ElectionDay #ElectionNight #Vote2016 #vote #USElection2016  https://t.
mlynne3||0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #ElectionDay #ElectionNight #Vote2016 #vote #USElection2016  https://t.
_saaaabs|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
_saaaabs|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
KellyFerg24|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
HelloTiffi_|ShopSeasonCaps|0.0|0.0|1.0|0.0|"RT @ShopSeasonCaps: Now Introducing the Red ""Hillary Blinton"" CapShop: https://t.co/EWOPpJ2hVb https://t.co/wjq7jULjyn"
HelloTiffi_|SeasonCaps|0.0|0.0|1.0|0.0|"RT @ShopSeasonCaps: Now Introducing the Red ""Hillary Blinton"" CapShop: https://t.co/EWOPpJ2hVb https://t.co/wjq7jULjyn"
michaelgmadden|romero|0.765|0.0|0.663|0.337|"RT @romero: If Hillary wins, I hope today will go down as Taco Tuesday. #HispanicVote #tacotuesday"
SMcCaulsky|humblethepoet|0.5719|0.0|0.709|0.291|RT @humblethepoet: If Hillary wins #Florida It's a wrap#electionday #ElectionNight #HERstory
berniebabe2016|mitchellvii|0.4404|0.0|0.861|0.139|RT @mitchellvii: I'm noticing the exit polls from MSNBC are dramatically better for Hillary than the ones from Fox.
holly_sebastian|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
holly_sebastian|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
lilla_ninni|jordanbrak|0.0268|0.3|0.433|0.267|"RT @jordanbrak: If Hillary wins I won't celebrate that she won, However I will celebrate that Trump lost #ElectionNight"
sn0wba111|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
ntvnyr173|mitchellvii|-0.7645|0.32|0.68|0.0|"RT @mitchellvii: Based upon exits, voters very unhappy with big money corruption.  That's bad for Hillary."
frazier_ann|newsbusters|0.8074|0.0|0.644|0.356|RT @newsbusters: Eleanor Clift Gushes Hillary Survived 'Hazing...With Stamina and Grace' On the Edge of Victory https://t.co/tNgTHDOOTP htt
frazier_ann|newsbusters|0.8074|0.0|0.644|0.356|RT @newsbusters: Eleanor Clift Gushes Hillary Survived 'Hazing...With Stamina and Grace' On the Edge of Victory https://t.co/tNgTHDOOTP htt
verdelishJP|boreanazs|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
verdelishJP|vine|-0.0191|0.097|0.903|0.0|RT @boreanazs: hillary and trump will never reach this level  https://t.co/H5WvbUT7ab
BrockGunn|TheOneandOnIyUS|0.7096|0.0|0.753|0.247|RT @TheOneandOnIyUS: The joke is on Hillary if she wins. She'll have to sit at the desk Monica sat under.
sliman12|StephensWSJ|0.8225|0.0|0.636|0.364|@StephensWSJ @WSJ Bret for the next 4 yrs you will have to justify your support of Hillary. Good luck.
DVader30|YoungDems4Trump|0.9042|0.0|0.621|0.379|"@YoungDems4Trump We wish Hillary well. If she wins, she wins. But the WHOLE Country will be watching each of her actions. Can she manage?"
grandmaj2|Pamela_Moore13|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
grandmaj2|twitter|0.0|0.0|1.0|0.0|RT @Pamela_Moore13: BREAKING:  Trump leads Hillary Clinton 52-41 in New Hampshire! https://t.co/dRUYoCaf3i
salberola|AFP|0.0|0.0|1.0|0.0|"RT @AFP: A large Hillary for America sign is displayed at the Jacob K. Javits Center in New York, where Clinton's #ElectionNight event is h"
frazman2|FuturisticHub|0.3436|0.151|0.616|0.233|@FuturisticHub @HillaryClinton Yeah. go ahead.. vote and loose.. Hillary fucked trump in his ass.. she is ma bitch.. :D D go hillary!!
johnscotthowell|YoungDems4Trump|0.2023|0.141|0.68|0.18|RT @YoungDems4Trump: if you are still undecided:Trump loves America.Hillary hates Americans.The choice is simple and clear.#myvote20
nickt1998|BroHumors|0.0|0.0|1.0|0.0|RT @BroHumors: Trump vs. Hillary  https://t.co/0jYBi7hlYO
nickt1998|vine|0.0|0.0|1.0|0.0|RT @BroHumors: Trump vs. Hillary  https://t.co/0jYBi7hlYO
saifuddinabd|mtredden|0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
saifuddinabd||0.0|0.0|1.0|0.0|"RT @mtredden: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https://"
vtoriac19|jordankerr23|0.8555|0.0|0.68|0.32|"RT @jordankerr23: Honestly though, how is Hillary supposed to take care of a country if she can't even take care of her teeth? https://t.co"
vtoriac19|t|0.8555|0.0|0.68|0.32|"RT @jordankerr23: Honestly though, how is Hillary supposed to take care of a country if she can't even take care of her teeth? https://t.co"
1kpook|XXL|0.34|0.0|0.821|0.179|RT @XXL: Kodak Black endorses Hillary Clinton from behind bars https://t.co/CnFMoKAN7M https://t.co/KPWegXMkdQ
1kpook|xxlmag|0.34|0.0|0.821|0.179|RT @XXL: Kodak Black endorses Hillary Clinton from behind bars https://t.co/CnFMoKAN7M https://t.co/KPWegXMkdQ
DaJourBrooks|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
tokiodaze|bawbbyspears|0.4404|0.0|0.674|0.326|RT @bawbbyspears: Hillary Clinton: *breathes*Trump supporters: https://t.co/UR1h1Gl9DM
tokiodaze|twitter|0.4404|0.0|0.674|0.326|RT @bawbbyspears: Hillary Clinton: *breathes*Trump supporters: https://t.co/UR1h1Gl9DM
SusanBugge|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
SusanBugge|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
JakeHober|PardonMyTake|0.5093|0.0|0.879|0.121|"RT @PardonMyTake: Hillary or Donald? Who cares, because In Canada we have all the chaw you could ever need. Come on over, America! We're so"
RadicalSamy|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
RadicalSamy|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
WackoTae313|imashbuttons|-0.0516|0.134|0.743|0.124|RT @imashbuttons: Why Hillary look like she bout to ask Yugi's grandpa bout some damn cards https://t.co/FZ4H3bLIoK
WackoTae313|twitter|-0.0516|0.134|0.743|0.124|RT @imashbuttons: Why Hillary look like she bout to ask Yugi's grandpa bout some damn cards https://t.co/FZ4H3bLIoK
WhosGoneGalt|BobMacAZ|0.2023|0.0|0.904|0.096|"RT @BobMacAZ: CIA Officially Breaks Their Silence, Reveals Top Secret Info on Hillary Shes Done https://t.co/oFQmT2ksXI via @USADailyInfo"
WhosGoneGalt|dailyinfo|0.2023|0.0|0.904|0.096|"RT @BobMacAZ: CIA Officially Breaks Their Silence, Reveals Top Secret Info on Hillary Shes Done https://t.co/oFQmT2ksXI via @USADailyInfo"
shadesofj0y|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
shadesofj0y|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
mvillz_|tylrmyrs|0.0|0.0|1.0|0.0|RT @tylrmyrs: Hillary on my paper ballotBernie on my heart ballot
808fong|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
808fong|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
mills_ann_julie|KGIRL0157|-0.5106|0.452|0.548|0.0|RT @KGIRL0157: Hillary for prison
EBChristyJr|TeamTrump|0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
EBChristyJr||0.6514|0.0|0.829|0.171|RT @TeamTrump: Hillary Clinton is simply unfit. It's time to put STRONG leadership in the White House - it's time to elect Trump!https://t
Duncaan17|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
squidninja|AMTrump4PRES|0.128|0.13|0.722|0.148|RT @AMTrump4PRES: #IAmVotingBecause My dad didn't sacrifice &amp; serve during 2 wars only 2C R great country become part of the #Hillary &amp; #So
YourstrulyBey|lilyachty|0.0|0.0|1.0|0.0|RT @lilyachty: Hillary! https://t.co/VZMLR24Y3Y
YourstrulyBey|twitter|0.0|0.0|1.0|0.0|RT @lilyachty: Hillary! https://t.co/VZMLR24Y3Y
niquuue|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
niquuue|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
Jennife40966102|JoyAnnReid|0.3182|0.0|0.887|0.113|RT @JoyAnnReid: Hillary Clinton being tied among white voters with a college degree is actually a huge swing toward Democrats. #ExitPolls
Jack2John|PhiKapMom|0.7603|0.0|0.783|0.217|RT @PhiKapMom: @AlGiordano Then you have the GOP women who won't tell their husband they voted for Hillary so great news!
bitchyologist|DanaSchwartzzz|0.6249|0.075|0.712|0.214|RT @DanaSchwartzzz: Dear lord if Hillary Clinton wins I'll read a book before bed and stop tweeting so much and give more to the homeless a
EastbTy|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
kamryn_hood|FemMajority|0.0|0.0|1.0|0.0|"RT @FemMajority: It's not just Hillary. Tonight, 7 women are trying to become the first female senator or house rep from their state: https"
goingscottyy|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
goingscottyy|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
vataormina|kmcwilliams5|0.7474|0.0|0.776|0.224|"RT @kmcwilliams5: And while you vote for Hillary Clinton explain to your future children why abortion at 36 weeks is legal, but not murder."
AshGotThis|mefeater|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
AshGotThis|twitter|0.5067|0.0|0.81|0.19|RT @mefeater: Big Freedia giving us a POLTICAL BOP! VOTE FOR HILLARY! VOTE FOR HILLARY! https://t.co/YwSS2vY5Xw
kentthonlo|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
ewwmeston|myboosartorius|0.0258|0.122|0.751|0.127|RT @myboosartorius: RT to be added into Hitlary's Hoes:-Must support Hillary Clinton-Talk about the election-No Dump Supporters-I'll be
juliacosta98|sofiercescotti|-0.2411|0.109|0.891|0.0|RT @sofiercescotti: im literally begging you if you havent votes yet please go vote Hillary i am afraid
rolaiamoda|DavidPapp|0.0|0.0|1.0|0.0|RT @DavidPapp: Photo of girl sleeping with Hillary Clinton action figure will melt your frozen heart https://t.co/tc0wWRMDCy
rolaiamoda|mashable|0.0|0.0|1.0|0.0|RT @DavidPapp: Photo of girl sleeping with Hillary Clinton action figure will melt your frozen heart https://t.co/tc0wWRMDCy
USAHipster|Koxinga8|0.7667|0.0|0.662|0.338|RT @Koxinga8: HAPPY ELECTION DAY! FBI Agents Just Surprised Comey With New Hillary Crimes https://t.co/Eafa46JVnq
USAHipster|angrypatriotmovement|0.7667|0.0|0.662|0.338|RT @Koxinga8: HAPPY ELECTION DAY! FBI Agents Just Surprised Comey With New Hillary Crimes https://t.co/Eafa46JVnq
lennnaaa_1|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
lennnaaa_1|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
JaviF7aca|rtsimpsons|0.0|0.0|1.0|0.0|RT @rtsimpsons: Ni Donald Trump ni Hillary Clinton. Lisa Simpson. https://t.co/COhFwMnSXq
JaviF7aca|twitter|0.0|0.0|1.0|0.0|RT @rtsimpsons: Ni Donald Trump ni Hillary Clinton. Lisa Simpson. https://t.co/COhFwMnSXq
WonderfulMaddie|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
WonderfulMaddie|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
tigersimon27|TIMENOUT|0.0|0.0|1.0|0.0|RT @TIMENOUT: WHY ARE ALL THE MACHINES SWITCHING TO HILLARY NOT TRUMP  Voters Reporting Ballots Switching To Clinton  https://t.co/nOm3v37
tigersimon27|t|0.0|0.0|1.0|0.0|RT @TIMENOUT: WHY ARE ALL THE MACHINES SWITCHING TO HILLARY NOT TRUMP  Voters Reporting Ballots Switching To Clinton  https://t.co/nOm3v37
RickVanWert|Stuboo3|0.0|0.0|1.0|0.0|@Stuboo3 Hillary Clinton eats Oreos without milk 
mprado1018|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
TrishFricke|LifeZette|0.4404|0.0|0.791|0.209|RT @LifeZette: Why @realDonaldTrump would be a better president for American women https://t.co/dyLBBgeB2c
TrishFricke|lifezette|0.4404|0.0|0.791|0.209|RT @LifeZette: Why @realDonaldTrump would be a better president for American women https://t.co/dyLBBgeB2c
DrThomasPaul|DrThomasPaul|0.6114|0.0|0.81|0.19|RT @DrThomasPaul: Happy about this #LGBT/#LGBTQ for anyone who thinks #Hillary is for #gays? Think again!She's financing #murders.#gayhttp
sydneylynnes|whytruy|-0.5106|0.113|0.887|0.0|RT @whytruy: vote hillary clinton idc if she a liar yall boyfriends lie to yall everyday &amp; yall still fw them so gone head &amp; vote for her
Halleywood|Dreamweasel|-0.7717|0.288|0.712|0.0|"RT @Dreamweasel: I predict they'll call it at 8:01 PST / 11:01 EST.Trump will concede defeat in about 5 years, and blame delay on Hillary"
SSNjl|linkis|-0.3382|0.138|0.862|0.0|"While Polls are Still Open, FBI Agents Drop the Biggest Bombshell Ever on HILLARY CLINTON! https://t.co/bpfEo4rzkN"
Raheemc_|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
eghofreshboi|tharealversace|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
eghofreshboi|twitter|0.0|0.0|1.0|0.0|RT @tharealversace: REASONS WHY YOU HAVE TO VOTE FOR HILLARY #VOTEHILLARY  https://t.co/eLzD2pVSw1
rachelkingmakeu|Lrihendry|0.7256|0.0|0.738|0.262|"RT @Lrihendry: Hillary supports this! If this is reason enough to support Trump, then you might want to sit this one out! #ElectionFina"
Cory21311812|nationdivided|-0.7959|0.336|0.664|0.0|RT @nationdivided: Indiana is joining Kentucky saying Hell No to Hillary! Go Trump #MAGA #Election2016 https://t.co/LvElXqBRef
Cory21311812|twitter|-0.7959|0.336|0.664|0.0|RT @nationdivided: Indiana is joining Kentucky saying Hell No to Hillary! Go Trump #MAGA #Election2016 https://t.co/LvElXqBRef
BGaideclin|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
BGaideclin|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
BreannaNicoleS8|AvesRyan|0.3612|0.0|0.848|0.152|RT @AvesRyan: Hillary Clinton becoming president is like Dan Scott becoming mayor of tree hill
guinnesssud|JaredWyand|-0.1027|0.057|0.943|0.0|RT @JaredWyand: The media wants to intimidate you into voting Hillary but nobody will know who you push that button forBreak the cycle #M
SusanNSunshine2|rollingstone|-0.0258|0.154|0.699|0.147|"Goes right along with hillary's ""cooking"".... no surprise.  #Freak  #ManBoobs  https://t.co/n7iI4eROSw https://t.co/YmrdZvuPUz"
unclebuckQPR|WillMcHoebag|0.3612|0.0|0.889|0.111|RT @WillMcHoebag: Hillary Clinton or Donald Trump? That's like asking whether you'd prefer Kate or Gerry McCann to babysit your kids.
sketjack|instagram|0.4724|0.0|0.796|0.204|Can't wait to see Hillary tonight!!!  Yall come join us at the https://t.co/Fb1dr0YVkd
Nikkie31479|AtlTeaPartyLove|0.0|0.0|1.0|0.0|"RT @AtlTeaPartyLove: If your Role Models are Jay Z, Beyonce and GaGa. You voted for Hillary because they told you to. Then, you already los"
bhola2063|Independent|0.0|0.0|1.0|0.0|RT @Independent: Where and when you can find the US presidential results https://t.co/VAMNBsX0VA
bhola2063|independent|0.0|0.0|1.0|0.0|RT @Independent: Where and when you can find the US presidential results https://t.co/VAMNBsX0VA
noahauten|memeprovider|-0.1695|0.196|0.804|0.0|"RT @memeprovider: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
boodaone1gmail1|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
boodaone1gmail1|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
Bhoysagoodin|CelticRockRoars|0.0|0.0|1.0|0.0|RT @CelticRockRoars: Woman on ITV just said people are blown away when they see Hillary.... everyone apart from Bill that is  #ElectionNig
sandysk53|INTJutsu|-0.5411|0.143|0.857|0.0|RT @INTJutsu: Hillary destroyed evidence after she received a subpoena to turn over all emails.  She should be in jail for that alone!#Ele
K_Ban|FelicityHuffman|0.7371|0.0|0.633|0.367|RT @FelicityHuffman: Voter loveWE LOVE HILLARY! @HillaryClinton #electionday #ImWithHer https://t.co/0AaJTaubSe
K_Ban|twitter|0.7371|0.0|0.633|0.367|RT @FelicityHuffman: Voter loveWE LOVE HILLARY! @HillaryClinton #electionday #ImWithHer https://t.co/0AaJTaubSe
Ian_Frado|_Coca_cole_a|0.5719|0.0|0.748|0.252|RT @_Coca_cole_a: If Hillary wins I'll give everyone who rt's this $5
joshua_economos|theScore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
joshua_economos|thescore|-0.5106|0.216|0.784|0.0|RT @theScore: Hornets' Spencer Hawes wears 'Hillary for Prison' shirt. #ElectionNight https://t.co/VYazSTvy4M https://t.co/mMq2j0bUig
andywtorre|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @ScottBaio @saskamare @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE NEW P
tragthagod|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
purplestar2015|FiveRights|-0.7783|0.274|0.726|0.0|"RT @FiveRights: #PodestaEmails35Hillary hates men, esp military men.Refused to meet w Lt Gen Sean MacFarland (top man in war against ISIS"
Feminismolizer|feminism|0.0|0.0|1.0|0.0|CNBC | Hillary Clinton 's unpopularity boils down to one... https://t.co/1WkIfk3dZk https://t.co/Skh2GXjW8I
_stylemuseum|twitter|0.0|0.0|1.0|0.0|Here&amp;rsquo;s How Kate McKinnon and Alec Baldwin Become Hillary Clinton and Donald Trump on Saturday https://t.co/8xanpkFQpW
KristiKotrous|KingsandLords|0.0|0.0|1.0|0.0|RT @KingsandLords: @MaddieAndMichi @enjoynChi @LilSteelerGirl @DebAlwaystrumpTRUMP 52%HillARY 43%JOHNSON 3%UNDECITED 2%USA LANDSLIDE
heeeeykidrauhl|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
Thatyguy955|FreddyAmazin|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
Thatyguy955|twitter|0.0|0.0|1.0|0.0|RT @FreddyAmazin: Rihanna wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  https://t.co/UFcFkP6js1
obe1cabo|qz|0.0|0.0|1.0|0.0|RT @qz: From Nina Simone to Beyonce: The Quartz playlist of songs by women who rule https://t.co/34y9D4BdxT
obe1cabo|qz|0.0|0.0|1.0|0.0|RT @qz: From Nina Simone to Beyonce: The Quartz playlist of songs by women who rule https://t.co/34y9D4BdxT
Da_La_Ca|Lexual__|0.3182|0.0|0.905|0.095|RT @Lexual__: Another comment: all the things y'all mentioned Hillary doing I'm sure Trump would have done if he had a career in politics.
irisheyes8701|mitchellvii|0.0|0.0|1.0|0.0|"RT @mitchellvii: Folks, in the two FL counties I've been watching, Hillary is DRAMATICALLY UNDERPERFORMING Obama.  We've got FL."
KimberlyFergus|JaredWyand|0.0|0.0|1.0|0.0|RT @JaredWyand: Hillary is on her way to an airport to watch the election results parked on a runway with flight plans to Qatar#ElectionD
TabataRouse|RedApplePol|0.5473|0.0|0.531|0.469|RT @RedApplePol: HERE'S HOPING  https://t.co/v0Yvnpt9hh
TabataRouse|aljazeera|0.5473|0.0|0.531|0.469|RT @RedApplePol: HERE'S HOPING  https://t.co/v0Yvnpt9hh
dianna_morales|ridevocals|-0.4588|0.146|0.778|0.075|"RT @ridevocals: WHY ARE PEOPLE VOTING TRUMP BECAUSE ""HILLARY IS A CRIMINAL"" WHEN THE FBI ALREADY CLEARED HER AND TRUMP IS GOING TO COURT FO"
alex_legue|ShuttupJenny|-0.1779|0.102|0.898|0.0|RT @ShuttupJenny: Rt if you keep having anxiety knowing Hillary Clinton might be elected president tomorrow
jayekasper|Sia|0.0|0.0|1.0|0.0|RT @Sia: VOTE FOR HILLARY #imwithher 
RhondaLorkowski|ChatRevolve|-0.296|0.091|0.909|0.0|RT @ChatRevolve: North Central I-4 Panhandle Tampa Tallahassee Florida get out and vote for Trump we need to stop Hillary Clinton | GO we n
F1Knox|DRUDGE_REPORT|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
F1Knox|businessinsider|0.0258|0.146|0.701|0.153|RT @DRUDGE_REPORT: VIDEO: CNN Reporter Shocked Female Voter Not Excited for Hillary... https://t.co/aZtk3j2TsN
Mari_Martinez08|Avstvn|-0.1695|0.196|0.804|0.0|"RT @Avstvn: We don't want Trump, we don't want Hillary, we just want Cory back in the house."
prepper1776|_HankRearden|0.2732|0.0|0.905|0.095|"RT @_HankRearden: I live in deep blue Boulder, in probably the bluest neighborhood. I've seen literally two Hillary signs total. The energy"
FergCapone|BangYaBrainsOut|0.5719|0.0|0.748|0.252|RT @BangYaBrainsOut: if Hillary wins I'll PayPal everyone $100 that RTs this.
xRomesMamax|TMITCH______|0.34|0.096|0.75|0.154|RT @TMITCH______: If Hillary wins she'll have to sit at the desk Monica sat under topping her man off smh
oxajc|TheHappyCampers|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
oxajc|twitter|0.8126|0.0|0.519|0.481|RT @TheHappyCampers: If Trump wins and if Hillary wins https://t.co/5HIZ9k3fZN
jrev2001|Whats_versace|0.5719|0.0|0.829|0.171|RT @Whats_versace: If Trump or Hillary  Wins The Election I Am Moving  Out Of The Country  Goodbye America  Hello   Uni
ejoy2270|Linnlondon1|-0.1111|0.117|0.783|0.101|RT @Linnlondon1: WARNING: MSM will call the election early in favor of Hillary to suppress Trump turnout. Don't listen. Get in line. Stay i
JLCole55|mitchellvii|0.5719|0.0|0.866|0.134|"RT @mitchellvii: Obama won FL by 73,000 votes in 2012.  So far, Hillary is behind Obama's 2012 pace by 60,000 votes IN JUST TWO COUNTIES. T"
imani_murray|RuffneckRefugee|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
imani_murray|t|-0.6486|0.163|0.837|0.0|RT @RuffneckRefugee: when trump will send you on the first boat back home but hillary will bomb you when you get there. https://t.co/rd3Sis
skylarariannaa|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
skylarariannaa|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
jiffyforthewin|MatthewKick|0.0|0.0|1.0|0.0|RT @MatthewKick: Choosing between Trump and Hillary #ElectionDay #myvote2016 https://t.co/JrPa4gKJBj
jiffyforthewin|twitter|0.0|0.0|1.0|0.0|RT @MatthewKick: Choosing between Trump and Hillary #ElectionDay #myvote2016 https://t.co/JrPa4gKJBj
Leo_eight20|infowars|-0.5719|0.346|0.654|0.0|RT @infowars: Even Kids Hate @HillaryClinton - https://t.co/X3GM45Gmjr #ElectionNight
Leo_eight20|infowars|-0.5719|0.346|0.654|0.0|RT @infowars: Even Kids Hate @HillaryClinton - https://t.co/X3GM45Gmjr #ElectionNight
EnjoiKimboh|ParksPics|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
EnjoiKimboh|twitter|0.0|0.0|1.0|0.0|RT @ParksPics: BREAKING HILLARY CLINTON NEWS THAT COULD COST HER THE ELECTION https://t.co/tdjwZ6McOc
estarr143|KaneZipperman|-0.6067|0.223|0.722|0.055|"RT @KaneZipperman: we don't care about Trump, we don't care about Hillary, we just want Cory back in the house"
matthew_sugg|maakaylakellyyy|0.0|0.0|1.0|0.0|RT @maakaylakellyyy: Voting for Hillary means... https://t.co/ziP1Q9RVrQ
matthew_sugg|twitter|0.0|0.0|1.0|0.0|RT @maakaylakellyyy: Voting for Hillary means... https://t.co/ziP1Q9RVrQ
Mystery77333|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
pmarcou3|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
pmarcou3|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
madirose_17|twitter|0.0|0.0|1.0|0.0|hillary #ImWithHer https://t.co/uf3XpC5WTy
calvinksbieber|Laughbook|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
calvinksbieber|twitter|-0.0191|0.089|0.911|0.0|RT @Laughbook: Trump and Hillary will never reach this level #electionday https://t.co/UqM6dObmZg
kim_means_gold|kim_means_gold|0.0|0.0|1.0|0.0|@kim_means_gold Way to go Hillary!
FuckBillyyyyyyy|chulomang|0.6207|0.0|0.78|0.22|RT @chulomang: Donald Trump Hillary Clinton Chief Keef DO YOU WANT REAL CHANGE? THERE IS A SOLUTION VOTE CHIEF KEEF #Election201
Sam_Giaccone|jess_rahth|-0.1263|0.181|0.667|0.152|RT @jess_rahth: Hillary looks like she'd be a really annoying and overly involved grandma
dmcveyy|KelseyKrause4|-0.1027|0.104|0.808|0.088|"RT @KelseyKrause4: if hillary was a male she would not be near as supported as she is, and that's the problem with modern feminism."
Svarela|TallahForTrump|-0.6229|0.338|0.662|0.0|RT @TallahForTrump: Don't vote for Hillary!She kills black people!#Haiti#BlackLivesMatter#ElectionDay#myvote2016
BobbyRuggles7|WSHHcomedy|0.0|0.0|1.0|0.0|RT @WSHHcomedy: Who's gonna be president? Hillary ??? LMAOOOOOOOO https://t.co/Q4SphHOiVS
BobbyRuggles7|twitter|0.0|0.0|1.0|0.0|RT @WSHHcomedy: Who's gonna be president? Hillary ??? LMAOOOOOOOO https://t.co/Q4SphHOiVS
IittIecurl|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
IittIecurl|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
davidpsdem|NelsyUmanzor|0.296|0.0|0.891|0.109|RT @NelsyUmanzor: Its #ElectionDay Join millions of Americans to vote for Hillary. Find out where you'll vote: https://t.co/b78xVeoTHl #Im
davidpsdem|iwillvote|0.296|0.0|0.891|0.109|RT @NelsyUmanzor: Its #ElectionDay Join millions of Americans to vote for Hillary. Find out where you'll vote: https://t.co/b78xVeoTHl #Im
nae3x_|novhak_|-0.6876|0.318|0.682|0.0|RT @novhak_: GO AWFFFFF Hillary !!!!!!! ( with your thick ass ) https://t.co/09fuQsvRaP
nae3x_|twitter|-0.6876|0.318|0.682|0.0|RT @novhak_: GO AWFFFFF Hillary !!!!!!! ( with your thick ass ) https://t.co/09fuQsvRaP
OldManDuke|Breaking911|-0.128|0.231|0.769|0.0|@Breaking911 Did #Hillary rig the election?
antonydeveaux|FrankLuntz|0.296|0.0|0.901|0.099|"RT @FrankLuntz: Michigan is going to end up for Hillary tonight.  I changed my opinion after seeing new numbers.Oh, and spoiler alert.  #"
savagecarlos___|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
savagecarlos___|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
Jennife30635376|AMTrump4PRES|0.128|0.13|0.722|0.148|RT @AMTrump4PRES: #IAmVotingBecause My dad didn't sacrifice &amp; serve during 2 wars only 2C R great country become part of the #Hillary &amp; #So
RUSTEAZY|souljaboy|-0.5719|0.493|0.19|0.318|RT @souljaboy: I hope Hillary win fuck trump stupid ass
aubnastyyy|EJKallenbach|0.0|0.0|1.0|0.0|RT @EJKallenbach: Imagine not having to hear about Hillary Clinton anymore  https://t.co/bfperX1jHQ
aubnastyyy|twitter|0.0|0.0|1.0|0.0|RT @EJKallenbach: Imagine not having to hear about Hillary Clinton anymore  https://t.co/bfperX1jHQ
JMemblatt|Caveman2743|0.4466|0.0|0.827|0.173|"RT @Caveman2743: RED ALERT: On Eve of Election, Benghazi BOMBSHELL Rains Down on Hillary https://t.co/rGox20vXgM"
JMemblatt|conservativetribune|0.4466|0.0|0.827|0.173|"RT @Caveman2743: RED ALERT: On Eve of Election, Benghazi BOMBSHELL Rains Down on Hillary https://t.co/rGox20vXgM"
jaleenmiller12|GIRLHEFUNNY|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
jaleenmiller12|twitter|-0.5106|0.202|0.798|0.0|RT @GIRLHEFUNNY: When they tell you don't vote for Hillary because she a liar  https://t.co/We2oiHoHy9
USAFMEDIC21|trump_florida|0.4019|0.0|0.828|0.172|RT @trump_florida: Source: The Military Times951 Active Duty Troops PolledTrump 54%     Hillary 25%#TrumpPence16 https://t.co/t1n374qx7M
USAFMEDIC21|twitter|0.4019|0.0|0.828|0.172|RT @trump_florida: Source: The Military Times951 Active Duty Troops PolledTrump 54%     Hillary 25%#TrumpPence16 https://t.co/t1n374qx7M
WyattMarsau|MattGallardo|-0.5859|0.352|0.648|0.0|RT @MattGallardo: Hillary Clinton will ruin our country.
dianebargar|HillaryClinton|-0.5267|0.268|0.732|0.0|"@HillaryClinton @mariobatali voted for Hillary, eating Mexican food, no wall No Trump.  Watching results"
studyequalmagic|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
johnvelasquez02|mariagross02|0.0772|0.0|0.874|0.126|@mariagross02 @cmmeyer221 obviously you want Hillary bc she's grandma too
smarquez58|WeLoveRobDyrdek|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
smarquez58|vine|0.0|0.0|1.0|0.0|RT @WeLoveRobDyrdek: When you have to vote for Trump or Hillary #ElectionDay https://t.co/khWIuhyETH
bopworldmag|zachhaller|-0.91|0.385|0.615|0.0|"RT @zachhaller: Blows my mind how many think the mean things Trump has saidare somehow worse than Hillary's career of lies, war, &amp; greed"
IDOLMADONNA|nytimes|0.7351|0.0|0.69|0.31|"RT @nytimes: Madonna played a surprise concert in New York last night, pledging her support for Hillary Clinton https://t.co/yHW261LrL1 htt"
IDOLMADONNA|nytimes|0.7351|0.0|0.69|0.31|"RT @nytimes: Madonna played a surprise concert in New York last night, pledging her support for Hillary Clinton https://t.co/yHW261LrL1 htt"
SamlCasper|rtsimpsons|0.0|0.0|1.0|0.0|RT @rtsimpsons: Ni Donald Trump ni Hillary Clinton. Lisa Simpson. https://t.co/COhFwMnSXq
SamlCasper|twitter|0.0|0.0|1.0|0.0|RT @rtsimpsons: Ni Donald Trump ni Hillary Clinton. Lisa Simpson. https://t.co/COhFwMnSXq
hrhpev|realAngeloGomez|0.25|0.0|0.778|0.222|@realAngeloGomez @monares_10 Hillary is endorsed by more fascists...https://t.co/SlPQR9bs0C
hrhpev|youtube|0.25|0.0|0.778|0.222|@realAngeloGomez @monares_10 Hillary is endorsed by more fascists...https://t.co/SlPQR9bs0C
DavidDeanLee1|2ALAW|-0.5859|0.192|0.808|0.0|RT @2ALAW: Voter Fraud In PhiladelphiaPush Button One For HillaryPaid For By The Democratic County.#ElectionNight #DonaldTrump https:/
DavidDeanLee1||-0.5859|0.192|0.808|0.0|RT @2ALAW: Voter Fraud In PhiladelphiaPush Button One For HillaryPaid For By The Democratic County.#ElectionNight #DonaldTrump https:/
randolphyuen731|satin_silkn|-0.2732|0.116|0.884|0.0|"RT @satin_silkn: While Polls Are Open, FBI Agents Drop The Biggest Bombshell Ever On Hillary Clinton https://t.co/1PdRYwjZZI"
randolphyuen731|redstatewatcher|-0.2732|0.116|0.884|0.0|"RT @satin_silkn: While Polls Are Open, FBI Agents Drop The Biggest Bombshell Ever On Hillary Clinton https://t.co/1PdRYwjZZI"
crustyJaureguii|TorisNormani|0.0|0.0|1.0|0.0|RT @TorisNormani: Either Trump or Hillary is gonna be president. U not voting isnt gonna change that. Even if only 1000 people voted it'd b
Asianpers_asion|RWF_10|0.4084|0.06|0.818|0.122|RT @RWF_10: It's one thing to SUPPORT Hillary over D. Trump. But to say &amp; believe she is not a corrupt &amp; manipulative human being seriously
AdorkableMazeau|twitter|0.7424|0.073|0.652|0.276|"A vote so profound, it brought three strangers to tears over the joy of voting for Hillary. I'm a proud democrat!  https://t.co/BpnLWA0Ss7"
DanielANestorJr|DontTread_2nd|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
DanielANestorJr|twitter|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
lopatonok|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
lopatonok|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
DanainFL|charliekirk11|-0.5255|0.34|0.486|0.175|RT @charliekirk11: RT if you proudly rejected the criminal that is Hillary Clinton!
becca_lynn|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
becca_lynn|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
ashleyroseeeee|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
ashleyroseeeee|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
kirstenadelmann|twitter|-0.3517|0.347|0.441|0.212|I don't like Hillary but this is funny as fuck HAHAHAHAHAHA https://t.co/oshYenwJGy
risejaeb|vickto_willy|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
risejaeb|t|-0.1531|0.109|0.806|0.085|"RT @vickto_willy: Hillary: ""Vote for me.""Me mimicking her: ""Vote for m- SHUT UP. You know damn well you the only option."" https://t.co/0OA"
Davietonner|DontTread_2nd|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
Davietonner|twitter|0.0|0.0|1.0|0.0|RT @DontTread_2nd: @Rambobiggs Is it connected to Hillary https://t.co/ruLA5yOK3k
September_Babe_|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
September_Babe_|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
FreedomTribe15|ed_hooley|0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #ElectionDay #ElectionNight #Vote2016 #vote #USElection2016  https://t.
FreedomTribe15||0.5267|0.0|0.761|0.239|RT @ed_hooley: Hillary Clinton &amp; John Podesta Spirit Cooking Party #ElectionDay #ElectionNight #Vote2016 #vote #USElection2016  https://t.
TwiloGuy73|0hour|0.2023|0.144|0.678|0.178|RT @0hour: Love how Twitter is reloading pro Hillary hashtags from months ago such losers in Silicon Valley.
ALEXswag97|J4CKMULL|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
ALEXswag97|twitter|0.0|0.0|1.0|0.0|RT @J4CKMULL: Hillary Clinton really did the #MannequinChallenge on #ElectionDay https://t.co/DxtJuf0zG0
MatKinman|youtube|0.0|0.0|1.0|0.0|Voting machines in Pennsylvania switch Trump votes to Hillary https://t.co/hyDnfSbTqo
Peggy7172|kincannon_show|-0.5849|0.296|0.704|0.0|RT @kincannon_show: This is very bad for Hillary --&gt; https://t.co/lv5ybXLiHZ
Peggy7172|twitter|-0.5849|0.296|0.704|0.0|RT @kincannon_show: This is very bad for Hillary --&gt; https://t.co/lv5ybXLiHZ
jetblackvheart|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
jetblackvheart|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
Ifubaraboye_|MrAyeDee|0.5859|0.099|0.586|0.315|"RT @MrAyeDee: Electoral irregularities everywhere. Dems are truly dedicated to getting Hillary elected,  no matter what... https://t.co/lm6"
Ifubaraboye_|t|0.5859|0.099|0.586|0.315|"RT @MrAyeDee: Electoral irregularities everywhere. Dems are truly dedicated to getting Hillary elected,  no matter what... https://t.co/lm6"
_Jaylaaa|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
_Jaylaaa|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
j_young62|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
ryantripp929|TheBardockObama|0.4215|0.0|0.781|0.219|RT @TheBardockObama: I had a nice election t shirt design butHillary Clinton deleted it.
BrandiBalls|CloydRivers|0.0|0.0|1.0|0.0|RT @CloydRivers: Im not against a woman bein President. Im just against that woman bein Hillary Clinton. Merica.
golfnovels|C_Tower|0.0|0.0|1.0|0.0|RT @C_Tower: WATCH  DO NOT VOTE Until Youve Seen THIS Hillary Video  She Wants It DELETED https://t.co/HSlobT8Z0E #Blacks4Trump #Grandpa
golfnovels|endingthefed|0.0|0.0|1.0|0.0|RT @C_Tower: WATCH  DO NOT VOTE Until Youve Seen THIS Hillary Video  She Wants It DELETED https://t.co/HSlobT8Z0E #Blacks4Trump #Grandpa
BTeboe|agreatercountry|-0.2481|0.135|0.767|0.099|"RT @agreatercountry: Lying MSM, for the last month is telling us the Latino support was surging for Hillary. CNN Poll shows NOT TRUE!http"
delanie_souders|BlaireHanks|-0.3612|0.136|0.798|0.066|RT @BlaireHanks: 2016:Attack of clowns Mourning of a gorilla for 7 monthsJuju on that beat Donald trump &amp; HillaryPeople pretending to
LuisMGuerra1|2ALAW|0.0|0.0|1.0|0.0|"RT @2ALAW: It's Over Folks!! NYPD Blows Whistle On #Hillary, Has Enough Evidence To Put Her Away For Life.@steph93065@SandraTXAS@AMTrum"
SallysNailz|facebook|0.6774|0.0|0.805|0.195|"LOL, so THIS lady VOTING next TO me GOES ""I JUST WANT TO VOTE FOR HILLARY &amp; GET THE PRESIDENT OUT OF THE WAY,... https://t.co/Jt9PxRJ4ox"
lltowing|FredZeppelin12|0.4404|0.0|0.884|0.116|"RT @FredZeppelin12: This needs to be RT'dHillary Clinton: ""We're Going to Take Things Away From You on Behalf of the Common Good"" http:"
chasewilber|tjNowak13|0.8737|0.0|0.678|0.322|RT @tjNowak13: TO ALL HILLARY SUPPORTERS: Don't waste your time going to vote. CNN says she has already won! RT to spread the word
Chimp999|cedric_persaud|-0.6289|0.256|0.744|0.0|"@cedric_persaud @JamieRJN @WayneDupreeShow SO, YOU AGREER WITH HILLARY THAT ALL AMERICANS ARE STUPID"
aubreyuss|Halezzzzzzzzzzz|-0.1027|0.069|0.931|0.0|RT @Halezzzzzzzzzzz: #Trump2016because Hillary doesn't deserve to be the first female president. Women have worked too hard to be represent
hallman_j|BrandonWeichert|0.0|0.0|1.0|0.0|RT @BrandonWeichert: @theIWP @SebGorka @realDonaldTrump @BoSnerdley @seanhannity @ericbolling  @AnnCoulter Voting 4 Hillary is a vote for p
jucerbone|antoniodelotero|0.6486|0.204|0.318|0.478|@antoniodelotero if Hillary wins cop haters win soo
k8koubz|RuariWould|0.1343|0.143|0.617|0.24|"@RuariWould I also hate this huge feminist surge for Hillary..surely you would want a competent person for the job, regardless of gender"
ShakiraShakira_|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
ShakiraShakira_|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
__NS__00|HillaryClinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
__NS__00|hillaryclinton|0.0|0.0|1.0|0.0|RT @HillaryClinton: Everything weve worked toward comes down to today. RT this if you're voting for Hillary: https://t.co/jfd3CXLD1s https
pabplanalp|maxkgom|0.4215|0.0|0.891|0.109|RT @maxkgom: ideally? hillary clinton and donald trump eat magic fortune cookies and wake up in each others' bodies and learn to see things
duncanmacmartin|PLTC_PastLives|0.0|0.0|1.0|0.0|RT @PLTC_PastLives: #NYT gave #HillaryClinton VETO POWER on all quotes (the paper confirms everything with #Hillary before printing it):ht
LNPurdie|mitchellvii|-0.1779|0.109|0.81|0.081|RT @mitchellvii: All of these early media predictions assume Hillary is getting all the Dem votes and ignoring Trumps advantage with Indies.
luckinubu|YoungDems4Trump|0.0|0.0|1.0|0.0|"RT @YoungDems4Trump: 207 Bernie voters for Trump in Arizona, folks! Counts as 414! Eat your heart out Hillary! I'm deflating your lies!#Yo"
ShaoIinTheDJ|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
ShaoIinTheDJ|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
p_inkd|rebel2187|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
p_inkd|twitter|0.0|0.0|1.0|0.0|RT @rebel2187: Donald and Hillary made an appearance in US Gov today  https://t.co/zOJflct4WM
barbaratien|Culture_Head|0.0|0.0|1.0|0.0|".@Culture_Head @kelleycalkins, we're bonded: #Sisterhood of the #voting #pantsuit #WearWhiteToVote https://t.co/qJfIw9YhCE @ESTBLSHMNT Rocks"
barbaratien|nytimes|0.0|0.0|1.0|0.0|".@Culture_Head @kelleycalkins, we're bonded: #Sisterhood of the #voting #pantsuit #WearWhiteToVote https://t.co/qJfIw9YhCE @ESTBLSHMNT Rocks"
PursuingMciver|tannermuro|-0.4588|0.158|0.842|0.0|RT @tannermuro: trump panicked and had to copy melania's ballot. now both are voting for hillary https://t.co/fiFO5tSrMh
PursuingMciver|twitter|-0.4588|0.158|0.842|0.0|RT @tannermuro: trump panicked and had to copy melania's ballot. now both are voting for hillary https://t.co/fiFO5tSrMh
MsPyatt|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
MsPyatt|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
stunnasingh|imchriskelly|0.5106|0.0|0.784|0.216|RT @imchriskelly: Imagine being as strong as Hillary Clinton. Literally. I cannot imagine that.
Janineleach6600|hitgirl2now|0.2732|0.0|0.9|0.1|"RT @hitgirl2now: Although Hillary is doing well with white, college educated women, this one voted 4 Trump.  I actually read the Wikileaks"
shelbyyyyleeann|memeprovider|-0.1695|0.196|0.804|0.0|"RT @memeprovider: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
matthew_tison|RonGorham|-0.9131|0.407|0.593|0.0|RT @RonGorham: @Conflicts @TrumpTrain09 @jimsciutto SMH this is Sirius!! We cannot let Hillary win ! This woman is the devil! https://t.co/
matthew_tison|t|-0.9131|0.407|0.593|0.0|RT @RonGorham: @Conflicts @TrumpTrain09 @jimsciutto SMH this is Sirius!! We cannot let Hillary win ! This woman is the devil! https://t.co/
jaydeyasemin|AJENews|0.5859|0.0|0.84|0.16|"RT @AJENews: Hillary Clinton gets most votes in Guam, a tiny island that has been predicting US election winner since 1980 https://t.co/SIq"
jaydeyasemin|t|0.5859|0.0|0.84|0.16|"RT @AJENews: Hillary Clinton gets most votes in Guam, a tiny island that has been predicting US election winner since 1980 https://t.co/SIq"
DrThomasPaul|DrThomasPaul|0.25|0.0|0.92|0.08|RT @DrThomasPaul: #Election2016 is the one where we set our differences aside and do the right thing. #Trump is the last chance for #Americ
golfnovels|newswirenet|-0.34|0.156|0.844|0.0|RT @newswirenet: Were the Iran Nuclear Negotiations Compromised by a Leak? https://t.co/1wB3eC0b7i #Hillary #Trump #Vote
golfnovels|newswire|-0.34|0.156|0.844|0.0|RT @newswirenet: Were the Iran Nuclear Negotiations Compromised by a Leak? https://t.co/1wB3eC0b7i #Hillary #Trump #Vote
ChampionNewsNet|cnn|0.0|0.0|1.0|0.0|My final 19 hours on the campaign trail with Clinton - https://t.co/PPgvSXwtHp
_paolamichele_|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
nicxdao|BuzzFeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
nicxdao|buzzfeed|0.0|0.0|1.0|0.0|RT @BuzzFeed: Rihanna just wore a shirt of herself wearing a Hillary Clinton shirt https://t.co/TFr2UJjW7n https://t.co/plOF0TDy1M
wiselatinaslink|twitter|0.4019|0.0|0.847|0.153|Hillary Clinton will treat women as equals. You know what Trump thinks of us. #ElectionNight https://t.co/jgMQt6sGbk
R666LEY|KayzoMusic|0.765|0.0|0.68|0.32|RT @KayzoMusic: If Hillary Clinton wins I hope she comes out for her victory speech to jotaro.
WasForBernie|WeAIIWin|0.0|0.0|1.0|0.0|"RT @WeAIIWin: @WWEAP25 Its @CNN, they @ananavarro provably work for the DNC/Hillary. Its Clinton News Network."
DiSwanson77|LibertyHacking|0.6208|0.084|0.671|0.245|RT @LibertyHacking: They're saying Trumps should respect the democratic system. SCREW THAT. Tell Hillary to respect the frigging law. #Elec
LeaningMike|twitter|0.0|0.0|1.0|0.0|"Hillarys own actions, obviously, had NOTHING to do with it.  What a sham.  CNN still spinning it. https://t.co/whNkfqZ0vn"
JR777771|hermanbutler1|0.2263|0.14|0.676|0.184|RT @hermanbutler1: Robert Reich: Dont Worry Hillary Clinton Will Win The Election https://t.co/hsSBwZoLUr #TNTweeters #USLatino #uniteblue
JR777771|linkis|0.2263|0.14|0.676|0.184|RT @hermanbutler1: Robert Reich: Dont Worry Hillary Clinton Will Win The Election https://t.co/hsSBwZoLUr #TNTweeters #USLatino #uniteblue
hebakhedr__|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
rebeca3436|Trapory|-0.8441|0.269|0.731|0.0|RT @Trapory: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
sandysk53|twitter|-0.7685|0.372|0.528|0.101|"Well, the way Hillary let 4 Americans die needlessly in BENGAZI REALLY BOTHERS ME! https://t.co/qmgl9ytOmb"
robison_gail|AlwayanAmerican|0.0|0.0|1.0|0.0|"RT @AlwayanAmerican: @IngrahamAngle @cubans4you Of Course not Obama , Hillary &amp; Voting Machines all belong to wanted Russian Fugitive Georg"
_WeLikeIke|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
_WeLikeIke|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
Katelynrossi3|kaleigh_ladner|-0.7003|0.281|0.667|0.052|"RT @kaleigh_ladner: No matter what happens today, I still hate Hillary Clinton, nothing will ever change my mind:)"
liquortroye|NeoXOver|0.8126|0.0|0.739|0.261|RT @NeoXOver: If Hillary wins I'll send Pizza Hut-promo codes to those who RTs this.If Trump wins I'll send Dominos-promo codes to those
david_macedo|DabneyPorte|-0.3818|0.126|0.874|0.0|RT @DabneyPorte: #ElectionNight #ExitPolls 45% who dislike both Trump and Hillary voted for TRUMP w only 27% choosing Hillary. WE A
Cr33perGal|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
lilliecorvs|Jamie_Daniels17|0.0772|0.0|0.843|0.157|"@Jamie_Daniels17 Hillary is a babe , rate her mannequin challenge "
Pedropjsn|rhm1947|-0.5574|0.247|0.753|0.0|"RT @rhm1947: Hillary Clinton ""We Came, We Saw, He Died"" (Gaddafi) https://t.co/whwiwbM22N"
Pedropjsn|linkis|-0.5574|0.247|0.753|0.0|"RT @rhm1947: Hillary Clinton ""We Came, We Saw, He Died"" (Gaddafi) https://t.co/whwiwbM22N"
societygirl123|USAMeg1|0.0|0.0|1.0|0.0|RT @USAMeg1: #FoxNews2016 Hillary Clinton belongs in jail not the Oval Office
WiredExGOP|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
tericento|AprilHayes_|-0.4724|0.139|0.861|0.0|RT @AprilHayes_: Stay in line West Coast!No to Hillary in the Primary! No in the General!#ElectionNight #Election2016 #iVoted #MAGAx3 #Ji
LennieJarratt|cnn|0.0|0.0|1.0|0.0|My final 19 hours on the campaign trail with Clinton https://t.co/22YlhsuInU
omezigue|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
omezigue|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
Azingra76|PrisonPlanet|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
Azingra76|twitter|-0.7251|0.303|0.697|0.0|RT @PrisonPlanet: More vote fraud in Philly. Dems handing out Hillary propaganda INSIDE polling station. https://t.co/CheWoAprKO
just_a_foody|FoxBusiness|0.5859|0.0|0.863|0.137|"RT @FoxBusiness: .@ktmcfarland: ""If [#Hillary] does win, she is not going to be able to govern. She has so much baggage, she is so corrupt."
Jacquel13895809|DrMartyFox|-0.5859|0.174|0.826|0.0|RT @DrMartyFox: #ImVotingBecause #Hillary Will Flood The Country With #Islamists Who Have Contempt For Our Culture #Christianity &amp; #Con
snouc|whytruy|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
snouc|twitter|0.3612|0.0|0.828|0.172|RT @whytruy: *casts vote for Hillary* Hillary: Thank you for your vot-Me: https://t.co/EjvxMWZD2c
MIACINO|justin_halpern|0.6476|0.0|0.751|0.249|RT @justin_halpern: My dream Hillary acceptance speech:*Bill introsBILL: The next president of the USA  (Borat voice) MA WIFE!HILLARY:
bvtgill|methwasp|0.5622|0.0|0.858|0.142|RT @methwasp: remember that a bill against abortion will only end SAFE abortions. remember that any reason you find to down hillary can be
Ianyb|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
SaraNaomie|broderick|0.6369|0.0|0.656|0.344|RT @broderick: Vine captured Hillary Clinton's best speech https://t.co/Iu0uyYheyz
SaraNaomie|vine|0.6369|0.0|0.656|0.344|RT @broderick: Vine captured Hillary Clinton's best speech https://t.co/Iu0uyYheyz
luckydbldd|JackPosobiec|-0.5574|0.265|0.735|0.0|RT @JackPosobiec: Illegal sign placement and Hillary worker placement everywhere https://t.co/pqrLmokcBn
luckydbldd|twitter|-0.5574|0.265|0.735|0.0|RT @JackPosobiec: Illegal sign placement and Hillary worker placement everywhere https://t.co/pqrLmokcBn
CARLOSIRUELA2|Pasion_Basket|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
CARLOSIRUELA2|twitter|0.0|0.0|1.0|0.0|"RT @Pasion_Basket: Ni Hillary Clinton, ni Donald Trump. JR SMITH FOR PRESIDENT!  https://t.co/0qhLtfR6wL"
ratstrash|urbandoll|0.0|0.0|1.0|0.0|@urbandoll didn't you previously say you were voting for Hillary or did i make this up in my head
Dnellzy|FunnyVines|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
Dnellzy|vine|-0.0191|0.089|0.911|0.0|RT @FunnyVines: Trump and Hillary will never reach this level #ElectionDay https://t.co/MqRHFPQCxh
yzzellmarieeee|memesuppIy|-0.1695|0.196|0.804|0.0|"RT @memesuppIy: We don't want Trump, we don't want Hillary, we just want Cory back in the house"
courtney_chid|The__Prototype|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
courtney_chid|twitter|-0.5719|0.236|0.764|0.0|RT @The__Prototype: Hillary: So y'all only with me cuz y'all hate Trump?Us: https://t.co/zqfFCAAOAV
BrianAmbler2|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
BrianAmbler2|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
maoamjetzt|jiujiuyulin|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
maoamjetzt|twitter|0.0516|0.154|0.679|0.167|RT @jiujiuyulin: The only convincing argument for Hillary I've heard all year. https://t.co/qGWJn3ygLt
ljarratt|cnn|0.0|0.0|1.0|0.0|My final 19 hours on the campaign trail with Clinton - https://t.co/J0k4RqHurn
ballerlife_7|_BeerPapi|0.8126|0.0|0.637|0.363|"RT @_BeerPapi: If Hillary wins, a bottle of henny.If Trump wins, a tall glass of bleach. https://t.co/VDVzCaZjvl"
ballerlife_7|twitter|0.8126|0.0|0.637|0.363|"RT @_BeerPapi: If Hillary wins, a bottle of henny.If Trump wins, a tall glass of bleach. https://t.co/VDVzCaZjvl"
manisterplan|PopCrave|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
manisterplan|twitter|0.0|0.0|1.0|0.0|RT @PopCrave: Rihanna wearing a shirt of her wearing a Hillary Clinton shirt is everything.  https://t.co/xqC3zfoJyZ
BeyonceMyRoc|twitter|0.6597|0.0|0.735|0.265|GA better have majorly voted for Hillary. I'm ready to pack my bags if they didn't https://t.co/Rz67cwxwQ6
Lilkimis1Legend|HoodBabyBop|-0.6211|0.177|0.752|0.072|RT @HoodBabyBop: #MyVote2016 is for my daughter who will know God and the kind of racist woman Hillary is!!! #VoteTrump I know Jesus is rea
snowm_|jacksfilms|0.8576|0.0|0.68|0.32|"RT @jacksfilms: ""If I win, I'm throwing you in jail!"" bellows Trump""Why?"" blushes Hillary""Because you're so sexy it's illegal""He then gr"
mayarajamani|twitter|0.0|0.0|1.0|0.0|"UES resident Jinji Nicole packed this jacket away years ago, but got it back out this year. ""It's my go-to fashion https://t.co/6ZBhPbJlJK"
casslyons24|twitter|0.0|0.0|1.0|0.0|A big (still bitter) F U to everyone that voted for Hillary instead of Bernie in the primaries  https://t.co/01zv6OysLi
JohnnyV213|Things4Guys|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
JohnnyV213|twitter|0.5719|0.0|0.761|0.239|RT @Things4Guys: Everyone's slamming Donald Trump but I didn't see Hillary Clinton help Kevin find the lobby https://t.co/mjZsOhLdhq
shivaputra|MODIvatingIndia|-0.6074|0.242|0.663|0.096|"RT @MODIvatingIndia: Dear, Trump &amp; Hillary, We don't care about you anymore. Our Prime Minister Modi dropped a NUCLEAR BOMB tonight. #Bla"
sam_govoni|JuiceTha56|0.168|0.0|0.927|0.073|RT @JuiceTha56: Will Hillary make pants suits mandatory? Will Trump build a wall on Mexicos border? Find out tomorrow on the season fin
alexfgravey|wikileaks|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
alexfgravey|regated|0.0|0.0|1.0|0.0|RT @wikileaks: Hillary Clinton is privately against gay marriage https://t.co/CvFM71cinV
Philly4Hillary|FrankLuntz|0.1571|0.091|0.792|0.117|RT @FrankLuntz: In case I wasn't clear enough from my previous tweets:Hillary Clinton will be the next President of the United States.  #
TyParkerS|shutupmikeginn|0.7227|0.0|0.771|0.229|@shutupmikeginn @GovGaryJohnson I think Hillary but maybe he'll come second in my precinct in la that's something to celebrate
rabbeni_kim|davidsirota|-0.2023|0.083|0.917|0.0|RT @davidsirota: Clinton Says She's Unaware Of Big Money That Oil And Gas Companies Have Given Her And Family Foundation https://t.co/xP27t
rabbeni_kim|t|-0.2023|0.083|0.917|0.0|RT @davidsirota: Clinton Says She's Unaware Of Big Money That Oil And Gas Companies Have Given Her And Family Foundation https://t.co/xP27t
elmerjfudd2012|Scarlett210|-0.765|0.28|0.72|0.0|"RT @Scarlett210: And #Hillary is a self-serving #elitist who'll continue #globalist policies, destroy ur safety&amp; deprive ur kids of a futur"
tezeqosycik|fentyy|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
tezeqosycik|twitter|0.0|0.0|1.0|0.0|RT @fentyy: Rihanna deadass wearing a t-shirt of herself wearing a t-shirt of Hillary Clinton  #ElectionDay https://t.co/OKngY7lvNs
ernierawlins2|GovMikeHuckabee|0.0|0.0|1.0|0.0|"RT @GovMikeHuckabee: State Dept says it takes 5 yrs to review 31,000 Hillary emails. Let Comey do it!  He can review 650,000 in 1 week!  ht"
messiah2kshow|nydailynews|0.3802|0.0|0.794|0.206|SEE IT! Madonna withdraws oral sex promise to Hillary voters  https://t.co/HG9AqnLwhm
StvnleyFlowers|LouisFarrakhan|0.2263|0.105|0.722|0.173|RT @LouisFarrakhan: You will find out that Hillary Clinton deceived you just like all of the rest before. They promise you everything and g
AnnaVi2001|philsadelphia|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
AnnaVi2001|twitter|0.7893|0.0|0.62|0.38|RT @philsadelphia: captain america voted for hillary so i think legally she should automatically win thank u https://t.co/cpkRZM1End
shivie|somhrd50|0.0|0.0|1.0|0.0|RT @somhrd50: I just told #NBCCT I voted today for Hillary #Clinton. Follow @nbcconnecticut for the latest election news.https://t.co/9izH
AriJameson|YoungDems4Trump|0.5994|0.0|0.824|0.176|RT @YoungDems4Trump: Dear Hillary voters on the fence. Think of our future. Think of her crimes against all of us. Please don't send us all
Boepperson|GreatAmericaPAC|0.0|0.0|1.0|0.0|RT @GreatAmericaPAC: Hear Dorothy Woods describe the stark difference between Trump and Crooked Hillary. https://t.co/biN5HhhpcO
Boepperson|twitter|0.0|0.0|1.0|0.0|RT @GreatAmericaPAC: Hear Dorothy Woods describe the stark difference between Trump and Crooked Hillary. https://t.co/biN5HhhpcO
tmmcgrath24|CloydRivers|-0.652|0.25|0.75|0.0|"RT @CloydRivers: Votin' for Hillary just because you don't like Trump, is like eatin' a turd just because you don't like broccoli. Merica."
rebecca_oyler|BandzUpDee|-0.8441|0.269|0.731|0.0|RT @BandzUpDee: Vote Hillary Clinton idc if she a liar y'all boyfriends lie to y'all everyday and y'all still fw them so VOTE HILLARY BITCH
Darksbane7|MamaJacquelyn|0.0|0.0|1.0|0.0|RT @MamaJacquelyn: Standing in line at 6:42am 7th person in line.  Can't wait to vote for Hillary!!!!!! #we'vegotthis
Zayshawn_Weston|AlexDonAudio|0.6739|0.0|0.807|0.193|RT @AlexDonAudio: WOW HILLARY JUST LOCKED IN THE BLACK VOTE FROM HALF COURT RT @RaeSremmurd: Go vote for her https://t.co/N8AHrXfpxV
Zayshawn_Weston|twitter|0.6739|0.0|0.807|0.193|RT @AlexDonAudio: WOW HILLARY JUST LOCKED IN THE BLACK VOTE FROM HALF COURT RT @RaeSremmurd: Go vote for her https://t.co/N8AHrXfpxV
ErikProgram|imashbuttons|-0.0516|0.134|0.743|0.124|RT @imashbuttons: Why Hillary look like she bout to ask Yugi's grandpa bout some damn cards https://t.co/FZ4H3bLIoK
ErikProgram|twitter|-0.0516|0.134|0.743|0.124|RT @imashbuttons: Why Hillary look like she bout to ask Yugi's grandpa bout some damn cards https://t.co/FZ4H3bLIoK
Colby_Howland|twitter|0.0|0.0|1.0|0.0|Who got into my phone?? It must had been Hillary.. #MakeAmericaGreatAgain #UpLikeDonaldTrump https://t.co/NtD0OJOJKK
